magic
tech scmos
timestamp 1731349415
<< nwell >>
rect 0 -6 25 26
<< ntransistor >>
rect 11 -22 13 -12
<< ptransistor >>
rect 11 0 13 20
<< ndiffusion >>
rect 6 -18 11 -12
rect 10 -22 11 -18
rect 13 -16 14 -12
rect 13 -22 18 -16
<< pdiffusion >>
rect 10 16 11 20
rect 6 0 11 16
rect 13 4 18 20
rect 13 0 14 4
<< ndcontact >>
rect 6 -22 10 -18
rect 14 -16 18 -12
<< pdcontact >>
rect 6 16 10 20
rect 14 0 18 4
<< polysilicon >>
rect 11 20 13 24
rect 11 -12 13 0
rect 11 -26 13 -22
<< polycontact >>
rect 7 -11 11 -7
<< metal1 >>
rect 0 27 25 30
rect 6 20 9 27
rect 15 -7 18 0
rect 0 -10 7 -7
rect 15 -10 22 -7
rect 15 -12 18 -10
rect 6 -27 9 -22
rect 0 -30 25 -27
<< labels >>
rlabel metal1 6 29 6 29 5 vdd
rlabel metal1 7 -29 7 -29 1 gnd
rlabel metal1 17 -8 17 -8 1 out
rlabel metal1 2 -9 2 -9 3 in
<< end >>
