.include TSMC_180nm.txt

.param SUPPLY=1.8
.global gnd vdd

VDD vdd gnd SUPPLY
vinA A gnd PULSE(0 SUPPLY   10ns 1ps 1ps   10ns  20ns)
vinB B gnd PULSE(0 SUPPLY    5ns 1ps 1ps    5ns  10ns)
vinC C gnd PULSE(0 SUPPLY  2.5ns 1ps 1ps  2.5ns   5ns)
vinD D gnd PULSE(0 SUPPLY 1.25ns 1ps 1ps 1.25ns 2.5ns)

.option scale=90n

M1000 gnd D a_1_n57# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=46u
M1001 vdd B output w_n28_n11# CMOSP w=20 l=2
+  ad=60p pd=26u as=60p ps=26u
M1002 vdd D output w_n28_n11# CMOSP w=20 l=2
+  ad=100p pd=50u as=60p ps=26u
M1003 output C vdd w_n28_n11# CMOSP w=20 l=2
+  ad=60p pd=26u as=60p ps=26u
M1004 output A vdd w_n28_n11# CMOSP w=20 l=2
+  ad=60p pd=26u as=100p ps=50u
M1005 a_n7_n57# B a_n15_n57# Gnd CMOSN w=40 l=2
+  ad=0.12n pd=46u as=0.12n ps=46u
M1006 a_1_n57# C a_n7_n57# Gnd CMOSN w=40 l=2
+  ad=0.12n pd=46u as=0.12n ps=46u
M1007 a_n15_n57# A output Gnd CMOSN w=40 l=2
+  ad=0.12n pd=46u as=0.2n ps=90u

.tran 1n 20n 

.control
  run
  set curplottitle="2024102023_4_NAND"
  * Plot output, and inputs shifted for visibility
  plot  v(A) v(B)+3 v(C)+6 v(D)+9 v(output)+12
.endc

.end