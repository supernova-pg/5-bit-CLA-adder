.include TSMC_180nm.txt

.param SUPPLY=1.8
.param LAMBDA=0.09u
.global gnd vdd

VDD vdd gnd SUPPLY
vinA A gnd PULSE(0 SUPPLY   20ns 1ps 1ps   20ns  40ns)
vinB B gnd PULSE(0 SUPPLY   10ns 1ps 1ps   10ns  20ns)
vinC C gnd PULSE(0 SUPPLY    5ns 1ps 1ps    5ns  10ns)
vinD D gnd PULSE(0 SUPPLY  2.5ns 1ps 1ps  2.5ns   5ns)
vinE E gnd PULSE(0 SUPPLY 1.25ns 1ps 1ps 1.25ns 2.5ns)

.option scale=90n

M1000 a_8_n73# C a_0_n73# gnd CMOSN w=50 l=2
+  ad=0.15n pd=56u as=0.15n ps=56u
M1001 a_n8_n73# A output gnd CMOSN w=50 l=2
+  ad=0.15n pd=56u as=0.25n ps=0.11m
M1002 a_16_n73# D a_8_n73# gnd CMOSN w=50 l=2
+  ad=0.15n pd=56u as=0.15n ps=56u
M1003 ground E a_16_n73# gnd CMOSN w=50 l=2
+  ad=0.25n pd=0.11m as=0.15n ps=56u
M1004 vdd D output w_n21_n15# CMOSP w=20 l=2
+  ad=60p pd=26u as=60p ps=26u
M1005 a_0_n73# B a_n8_n73# gnd CMOSN w=50 l=2
+  ad=0.15n pd=56u as=0.15n ps=56u
M1006 output A vdd w_n21_n15# CMOSP w=20 l=2
+  ad=60p pd=26u as=100p ps=50u
M1007 output C vdd w_n21_n15# CMOSP w=20 l=2
+  ad=60p pd=26u as=60p ps=26u
M1008 output E vdd w_n21_n15# CMOSP w=20 l=2
+  ad=100p pd=50u as=60p ps=26u
M1009 vdd B output w_n21_n15# CMOSP w=20 l=2
+  ad=60p pd=26u as=60p ps=26u



.tran 1n 80n 


.control

    run
    set curplottitle="2024102023_5_nand"
    plot v(A) v(B)+3 v(C)+6 v(D)+9 v(E)+12 v(output)+15
    
.endc
.end