magic
tech scmos
timestamp 1763554598
<< nwell >>
rect -21 -15 35 17
<< ntransistor >>
rect -10 -73 -8 -23
rect -2 -73 0 -23
rect 6 -73 8 -23
rect 14 -73 16 -23
rect 22 -73 24 -23
<< ptransistor >>
rect -10 -9 -8 11
rect -2 -9 0 11
rect 6 -9 8 11
rect 14 -9 16 11
rect 22 -9 24 11
<< ndiffusion >>
rect -11 -73 -10 -23
rect -8 -73 -7 -23
rect -3 -73 -2 -23
rect 0 -73 1 -23
rect 5 -73 6 -23
rect 8 -73 9 -23
rect 13 -73 14 -23
rect 16 -73 17 -23
rect 21 -73 22 -23
rect 24 -73 25 -23
<< pdiffusion >>
rect -11 -9 -10 11
rect -8 -9 -7 11
rect -3 -9 -2 11
rect 0 -9 1 11
rect 5 -9 6 11
rect 8 -9 9 11
rect 13 -9 14 11
rect 16 -9 17 11
rect 21 -9 22 11
rect 24 -9 25 11
<< ndcontact >>
rect -15 -73 -11 -23
rect -7 -73 -3 -23
rect 1 -73 5 -23
rect 9 -73 13 -23
rect 17 -73 21 -23
rect 25 -73 29 -23
<< pdcontact >>
rect -15 -9 -11 11
rect -7 -9 -3 11
rect 1 -9 5 11
rect 9 -9 13 11
rect 17 -9 21 11
rect 25 -9 29 11
<< polysilicon >>
rect -10 11 -8 14
rect -2 11 0 14
rect 6 11 8 14
rect 14 11 16 14
rect 22 11 24 14
rect -10 -23 -8 -9
rect -2 -23 0 -9
rect 6 -23 8 -9
rect 14 -23 16 -9
rect 22 -23 24 -9
rect -10 -81 -8 -73
rect -2 -81 0 -73
rect 6 -81 8 -73
rect 14 -81 16 -73
rect 22 -81 24 -73
<< polycontact >>
rect -11 -85 -7 -81
rect -3 -85 1 -81
rect 5 -85 9 -81
rect 13 -85 17 -81
rect 21 -85 25 -81
<< metal1 >>
rect -15 11 -11 13
rect 1 11 5 13
rect 17 11 21 13
rect -7 -10 -3 -9
rect 9 -10 13 -9
rect 25 -10 29 -9
rect -15 -23 -11 -21
rect 25 -74 29 -73
rect 25 -78 34 -74
rect -12 -90 -7 -85
rect -4 -90 1 -85
rect 4 -90 9 -85
rect 13 -90 18 -85
rect 21 -90 26 -85
<< m2contact >>
rect -15 13 -10 18
rect 1 13 6 18
rect 17 13 22 18
rect -7 -15 -2 -10
rect 9 -15 14 -10
rect 25 -15 30 -10
rect -16 -21 -11 -16
<< metal2 >>
rect -15 18 -11 27
rect -10 13 1 17
rect 6 13 17 17
rect -2 -15 9 -11
rect 14 -15 25 -11
rect -7 -16 -3 -15
rect -21 -20 -16 -16
rect -11 -20 -3 -16
<< labels >>
rlabel metal1 -12 -90 -7 -85 1 input_1
rlabel metal1 -4 -90 1 -85 1 input_2
rlabel metal1 4 -90 9 -85 1 input_3
rlabel metal1 13 -90 18 -85 1 input_4
rlabel metal1 21 -90 26 -85 1 input_5
rlabel metal1 29 -78 34 -74 7 ground
rlabel metal2 -21 -20 -16 -16 3 output
rlabel metal2 -15 18 -11 27 5 power
<< end >>
