magic
tech scmos
timestamp 1764710698
<< nwell >>
rect 38 957 70 1018
rect 17 896 49 928
rect 914 892 946 948
rect 43 859 75 884
rect 895 805 927 853
rect 38 741 70 802
rect 885 718 917 758
rect 1209 753 1241 809
rect 1649 737 1681 798
rect 17 680 49 712
rect 43 643 75 668
rect 850 652 882 684
rect 38 525 70 586
rect 897 540 929 588
rect 17 464 49 496
rect 887 463 919 503
rect 1203 459 1235 507
rect 43 427 75 452
rect 1641 437 1673 498
rect 850 400 882 432
rect 38 309 70 370
rect 888 300 920 340
rect 1205 285 1237 325
rect 1641 287 1673 348
rect 17 248 49 280
rect 851 237 883 269
rect 43 211 75 236
rect 849 154 881 186
rect 38 93 70 154
rect 1165 153 1197 185
rect 1641 149 1673 210
rect 17 32 49 64
rect 43 -5 75 20
<< ntransistor >>
rect 22 1005 32 1007
rect 21 977 31 979
rect 21 968 31 970
rect 856 935 906 937
rect 856 927 906 929
rect 856 919 906 921
rect 57 915 77 917
rect 856 911 906 913
rect 57 907 77 909
rect 856 903 906 905
rect 27 871 37 873
rect 849 840 889 842
rect 849 832 889 834
rect 849 824 889 826
rect 849 816 889 818
rect 1151 796 1201 798
rect 22 789 32 791
rect 1151 788 1201 790
rect 1633 785 1643 787
rect 1151 780 1201 782
rect 1151 772 1201 774
rect 1151 764 1201 766
rect 21 761 31 763
rect 1632 757 1642 759
rect 21 752 31 754
rect 1632 748 1642 750
rect 844 745 874 747
rect 844 737 874 739
rect 844 729 874 731
rect 57 699 77 701
rect 57 691 77 693
rect 890 671 910 673
rect 890 663 910 665
rect 27 655 37 657
rect 22 573 32 575
rect 851 575 891 577
rect 851 567 891 569
rect 851 559 891 561
rect 851 551 891 553
rect 21 545 31 547
rect 21 536 31 538
rect 1157 494 1197 496
rect 846 490 876 492
rect 57 483 77 485
rect 1157 486 1197 488
rect 846 482 876 484
rect 57 475 77 477
rect 846 474 876 476
rect 1625 485 1635 487
rect 1157 478 1197 480
rect 1157 470 1197 472
rect 1624 457 1634 459
rect 1624 448 1634 450
rect 27 439 37 441
rect 890 419 910 421
rect 890 411 910 413
rect 22 357 32 359
rect 1625 335 1635 337
rect 21 329 31 331
rect 847 327 877 329
rect 21 320 31 322
rect 847 319 877 321
rect 847 311 877 313
rect 1164 312 1194 314
rect 1624 307 1634 309
rect 1164 304 1194 306
rect 1624 298 1634 300
rect 1164 296 1194 298
rect 57 267 77 269
rect 57 259 77 261
rect 891 256 911 258
rect 891 248 911 250
rect 27 223 37 225
rect 1625 197 1635 199
rect 889 173 909 175
rect 1205 172 1225 174
rect 889 165 909 167
rect 1624 169 1634 171
rect 1205 164 1225 166
rect 1624 160 1634 162
rect 22 141 32 143
rect 21 113 31 115
rect 21 104 31 106
rect 57 51 77 53
rect 57 43 77 45
rect 27 7 37 9
<< ptransistor >>
rect 44 1005 64 1007
rect 44 977 64 979
rect 44 968 64 970
rect 920 935 940 937
rect 920 927 940 929
rect 920 919 940 921
rect 23 915 43 917
rect 920 911 940 913
rect 23 907 43 909
rect 920 903 940 905
rect 49 871 69 873
rect 901 840 921 842
rect 901 832 921 834
rect 901 824 921 826
rect 901 816 921 818
rect 1215 796 1235 798
rect 44 789 64 791
rect 1215 788 1235 790
rect 1655 785 1675 787
rect 1215 780 1235 782
rect 1215 772 1235 774
rect 1215 764 1235 766
rect 44 761 64 763
rect 1655 757 1675 759
rect 44 752 64 754
rect 1655 748 1675 750
rect 891 745 911 747
rect 891 737 911 739
rect 891 729 911 731
rect 23 699 43 701
rect 23 691 43 693
rect 856 671 876 673
rect 856 663 876 665
rect 49 655 69 657
rect 44 573 64 575
rect 903 575 923 577
rect 903 567 923 569
rect 903 559 923 561
rect 903 551 923 553
rect 44 545 64 547
rect 44 536 64 538
rect 1209 494 1229 496
rect 893 490 913 492
rect 23 483 43 485
rect 1209 486 1229 488
rect 893 482 913 484
rect 23 475 43 477
rect 893 474 913 476
rect 1647 485 1667 487
rect 1209 478 1229 480
rect 1209 470 1229 472
rect 1647 457 1667 459
rect 1647 448 1667 450
rect 49 439 69 441
rect 856 419 876 421
rect 856 411 876 413
rect 44 357 64 359
rect 1647 335 1667 337
rect 44 329 64 331
rect 894 327 914 329
rect 44 320 64 322
rect 894 319 914 321
rect 894 311 914 313
rect 1211 312 1231 314
rect 1647 307 1667 309
rect 1211 304 1231 306
rect 1647 298 1667 300
rect 1211 296 1231 298
rect 23 267 43 269
rect 23 259 43 261
rect 857 256 877 258
rect 857 248 877 250
rect 49 223 69 225
rect 1647 197 1667 199
rect 855 173 875 175
rect 1171 172 1191 174
rect 855 165 875 167
rect 1647 169 1667 171
rect 1171 164 1191 166
rect 1647 160 1667 162
rect 44 141 64 143
rect 44 113 64 115
rect 44 104 64 106
rect 23 51 43 53
rect 23 43 43 45
rect 49 7 69 9
<< ndiffusion >>
rect 26 1008 32 1012
rect 22 1007 32 1008
rect 22 1004 32 1005
rect 26 1000 32 1004
rect 25 980 31 984
rect 21 979 31 980
rect 21 976 31 977
rect 21 972 27 976
rect 21 970 31 972
rect 21 967 31 968
rect 21 963 27 967
rect 856 937 906 938
rect 856 934 906 935
rect 856 929 906 930
rect 856 926 906 927
rect 856 921 906 922
rect 856 918 906 919
rect 57 917 77 918
rect 57 914 77 915
rect 856 913 906 914
rect 856 910 906 911
rect 57 909 77 910
rect 57 906 77 907
rect 856 905 906 906
rect 856 902 906 903
rect 31 874 37 878
rect 27 873 37 874
rect 27 870 37 871
rect 27 866 33 870
rect 849 842 889 843
rect 849 839 889 840
rect 849 834 889 835
rect 849 831 889 832
rect 849 826 889 827
rect 849 823 889 824
rect 849 818 889 819
rect 849 815 889 816
rect 26 792 32 796
rect 22 791 32 792
rect 1151 798 1201 799
rect 1151 795 1201 796
rect 22 788 32 789
rect 26 784 32 788
rect 1151 790 1201 791
rect 1637 788 1643 792
rect 1151 787 1201 788
rect 1151 782 1201 783
rect 1633 787 1643 788
rect 1633 784 1643 785
rect 1637 780 1643 784
rect 1151 779 1201 780
rect 1151 774 1201 775
rect 1151 771 1201 772
rect 25 764 31 768
rect 21 763 31 764
rect 1151 766 1201 767
rect 1151 763 1201 764
rect 21 760 31 761
rect 21 756 27 760
rect 21 754 31 756
rect 1636 760 1642 764
rect 1632 759 1642 760
rect 1632 756 1642 757
rect 21 751 31 752
rect 21 747 27 751
rect 844 747 874 748
rect 1632 752 1638 756
rect 1632 750 1642 752
rect 1632 747 1642 748
rect 844 744 874 745
rect 844 739 874 740
rect 1632 743 1638 747
rect 844 736 874 737
rect 844 731 874 732
rect 844 728 874 729
rect 57 701 77 702
rect 57 698 77 699
rect 57 693 77 694
rect 57 690 77 691
rect 890 673 910 674
rect 890 670 910 671
rect 890 665 910 666
rect 31 658 37 662
rect 27 657 37 658
rect 890 662 910 663
rect 27 654 37 655
rect 27 650 33 654
rect 26 576 32 580
rect 22 575 32 576
rect 851 577 891 578
rect 851 574 891 575
rect 22 572 32 573
rect 26 568 32 572
rect 851 569 891 570
rect 851 566 891 567
rect 851 561 891 562
rect 851 558 891 559
rect 25 548 31 552
rect 21 547 31 548
rect 851 553 891 554
rect 851 550 891 551
rect 21 544 31 545
rect 21 540 27 544
rect 21 538 31 540
rect 21 535 31 536
rect 21 531 27 535
rect 846 492 876 493
rect 1157 496 1197 497
rect 1157 493 1197 494
rect 846 489 876 490
rect 57 485 77 486
rect 57 482 77 483
rect 846 484 876 485
rect 1157 488 1197 489
rect 1629 488 1635 492
rect 1625 487 1635 488
rect 1157 485 1197 486
rect 846 481 876 482
rect 57 477 77 478
rect 57 474 77 475
rect 846 476 876 477
rect 846 473 876 474
rect 1157 480 1197 481
rect 1625 484 1635 485
rect 1629 480 1635 484
rect 1157 477 1197 478
rect 1157 472 1197 473
rect 1157 469 1197 470
rect 1628 460 1634 464
rect 1624 459 1634 460
rect 1624 456 1634 457
rect 1624 452 1630 456
rect 1624 450 1634 452
rect 1624 447 1634 448
rect 31 442 37 446
rect 27 441 37 442
rect 1624 443 1630 447
rect 27 438 37 439
rect 27 434 33 438
rect 890 421 910 422
rect 890 418 910 419
rect 890 413 910 414
rect 890 410 910 411
rect 26 360 32 364
rect 22 359 32 360
rect 22 356 32 357
rect 26 352 32 356
rect 1629 338 1635 342
rect 1625 337 1635 338
rect 25 332 31 336
rect 21 331 31 332
rect 1625 334 1635 335
rect 21 328 31 329
rect 21 324 27 328
rect 21 322 31 324
rect 847 329 877 330
rect 1629 330 1635 334
rect 847 326 877 327
rect 21 319 31 320
rect 21 315 27 319
rect 847 321 877 322
rect 847 318 877 319
rect 847 313 877 314
rect 1164 314 1194 315
rect 1164 311 1194 312
rect 847 310 877 311
rect 1164 306 1194 307
rect 1628 310 1634 314
rect 1624 309 1634 310
rect 1624 306 1634 307
rect 1164 303 1194 304
rect 1164 298 1194 299
rect 1624 302 1630 306
rect 1624 300 1634 302
rect 1624 297 1634 298
rect 1164 295 1194 296
rect 1624 293 1630 297
rect 57 269 77 270
rect 57 266 77 267
rect 57 261 77 262
rect 57 258 77 259
rect 891 258 911 259
rect 891 255 911 256
rect 891 250 911 251
rect 891 247 911 248
rect 31 226 37 230
rect 27 225 37 226
rect 27 222 37 223
rect 27 218 33 222
rect 1629 200 1635 204
rect 1625 199 1635 200
rect 1625 196 1635 197
rect 1629 192 1635 196
rect 889 175 909 176
rect 889 172 909 173
rect 1205 174 1225 175
rect 1628 172 1634 176
rect 889 167 909 168
rect 889 164 909 165
rect 1205 171 1225 172
rect 1624 171 1634 172
rect 1205 166 1225 167
rect 1624 168 1634 169
rect 1205 163 1225 164
rect 1624 164 1630 168
rect 1624 162 1634 164
rect 1624 159 1634 160
rect 1624 155 1630 159
rect 26 144 32 148
rect 22 143 32 144
rect 22 140 32 141
rect 26 136 32 140
rect 25 116 31 120
rect 21 115 31 116
rect 21 112 31 113
rect 21 108 27 112
rect 21 106 31 108
rect 21 103 31 104
rect 21 99 27 103
rect 57 53 77 54
rect 57 50 77 51
rect 57 45 77 46
rect 57 42 77 43
rect 31 10 37 14
rect 27 9 37 10
rect 27 6 37 7
rect 27 2 33 6
<< pdiffusion >>
rect 48 1008 64 1012
rect 44 1007 64 1008
rect 44 1004 64 1005
rect 44 1000 60 1004
rect 44 980 60 984
rect 44 979 64 980
rect 44 976 64 977
rect 44 972 46 976
rect 50 972 64 976
rect 44 970 64 972
rect 44 967 64 968
rect 48 963 64 967
rect 920 937 940 938
rect 920 934 940 935
rect 920 929 940 930
rect 23 917 43 918
rect 920 926 940 927
rect 920 921 940 922
rect 23 914 43 915
rect 23 909 43 910
rect 920 918 940 919
rect 920 913 940 914
rect 23 906 43 907
rect 920 910 940 911
rect 920 905 940 906
rect 920 902 940 903
rect 49 874 65 878
rect 49 873 69 874
rect 49 870 69 871
rect 53 866 69 870
rect 901 842 921 843
rect 901 839 921 840
rect 901 834 921 835
rect 901 831 921 832
rect 901 826 921 827
rect 901 823 921 824
rect 901 818 921 819
rect 901 815 921 816
rect 48 792 64 796
rect 1215 798 1235 799
rect 44 791 64 792
rect 44 788 64 789
rect 44 784 60 788
rect 1215 795 1235 796
rect 1215 790 1235 791
rect 1215 787 1235 788
rect 1659 788 1675 792
rect 1655 787 1675 788
rect 1215 782 1235 783
rect 1655 784 1675 785
rect 1655 780 1671 784
rect 1215 779 1235 780
rect 1215 774 1235 775
rect 44 764 60 768
rect 44 763 64 764
rect 1215 771 1235 772
rect 1215 766 1235 767
rect 44 760 64 761
rect 44 756 46 760
rect 50 756 64 760
rect 1215 763 1235 764
rect 1655 760 1671 764
rect 1655 759 1675 760
rect 44 754 64 756
rect 44 751 64 752
rect 48 747 64 751
rect 1655 756 1675 757
rect 1655 752 1657 756
rect 1661 752 1675 756
rect 1655 750 1675 752
rect 891 747 911 748
rect 891 744 911 745
rect 1655 747 1675 748
rect 1659 743 1675 747
rect 891 739 911 740
rect 891 736 911 737
rect 891 731 911 732
rect 891 728 911 729
rect 23 701 43 702
rect 23 698 43 699
rect 23 693 43 694
rect 23 690 43 691
rect 856 673 876 674
rect 856 670 876 671
rect 856 665 876 666
rect 856 662 876 663
rect 49 658 65 662
rect 49 657 69 658
rect 49 654 69 655
rect 53 650 69 654
rect 48 576 64 580
rect 44 575 64 576
rect 903 577 923 578
rect 44 572 64 573
rect 44 568 60 572
rect 903 574 923 575
rect 903 569 923 570
rect 903 566 923 567
rect 903 561 923 562
rect 44 548 60 552
rect 903 558 923 559
rect 903 553 923 554
rect 44 547 64 548
rect 903 550 923 551
rect 44 544 64 545
rect 44 540 46 544
rect 50 540 64 544
rect 44 538 64 540
rect 44 535 64 536
rect 48 531 64 535
rect 23 485 43 486
rect 1209 496 1229 497
rect 893 492 913 493
rect 23 482 43 483
rect 23 477 43 478
rect 893 489 913 490
rect 1209 493 1229 494
rect 1209 488 1229 489
rect 1651 488 1667 492
rect 1647 487 1667 488
rect 893 484 913 485
rect 23 474 43 475
rect 893 481 913 482
rect 893 476 913 477
rect 893 473 913 474
rect 1209 485 1229 486
rect 1209 480 1229 481
rect 1647 484 1667 485
rect 1647 480 1663 484
rect 1209 477 1229 478
rect 1209 472 1229 473
rect 1209 469 1229 470
rect 1647 460 1663 464
rect 1647 459 1667 460
rect 1647 456 1667 457
rect 1647 452 1649 456
rect 1653 452 1667 456
rect 1647 450 1667 452
rect 49 442 65 446
rect 1647 447 1667 448
rect 1651 443 1667 447
rect 49 441 69 442
rect 49 438 69 439
rect 53 434 69 438
rect 856 421 876 422
rect 856 418 876 419
rect 856 413 876 414
rect 856 410 876 411
rect 48 360 64 364
rect 44 359 64 360
rect 44 356 64 357
rect 44 352 60 356
rect 1651 338 1667 342
rect 1647 337 1667 338
rect 44 332 60 336
rect 44 331 64 332
rect 44 328 64 329
rect 44 324 46 328
rect 50 324 64 328
rect 1647 334 1667 335
rect 1647 330 1663 334
rect 894 329 914 330
rect 44 322 64 324
rect 44 319 64 320
rect 48 315 64 319
rect 894 326 914 327
rect 894 321 914 322
rect 894 318 914 319
rect 894 313 914 314
rect 1211 314 1231 315
rect 894 310 914 311
rect 1211 311 1231 312
rect 1647 310 1663 314
rect 1647 309 1667 310
rect 1211 306 1231 307
rect 1211 303 1231 304
rect 1211 298 1231 299
rect 1647 306 1667 307
rect 1647 302 1649 306
rect 1653 302 1667 306
rect 1647 300 1667 302
rect 1211 295 1231 296
rect 1647 297 1667 298
rect 1651 293 1667 297
rect 23 269 43 270
rect 23 266 43 267
rect 23 261 43 262
rect 23 258 43 259
rect 857 258 877 259
rect 857 255 877 256
rect 857 250 877 251
rect 857 247 877 248
rect 49 226 65 230
rect 49 225 69 226
rect 49 222 69 223
rect 53 218 69 222
rect 1651 200 1667 204
rect 1647 199 1667 200
rect 1647 196 1667 197
rect 1647 192 1663 196
rect 855 175 875 176
rect 855 172 875 173
rect 855 167 875 168
rect 1171 174 1191 175
rect 1171 171 1191 172
rect 855 164 875 165
rect 1171 166 1191 167
rect 1647 172 1663 176
rect 1647 171 1667 172
rect 1171 163 1191 164
rect 1647 168 1667 169
rect 1647 164 1649 168
rect 1653 164 1667 168
rect 1647 162 1667 164
rect 1647 159 1667 160
rect 1651 155 1667 159
rect 48 144 64 148
rect 44 143 64 144
rect 44 140 64 141
rect 44 136 60 140
rect 44 116 60 120
rect 44 115 64 116
rect 44 112 64 113
rect 44 108 46 112
rect 50 108 64 112
rect 44 106 64 108
rect 44 103 64 104
rect 48 99 64 103
rect 23 53 43 54
rect 23 50 43 51
rect 23 45 43 46
rect 23 42 43 43
rect 49 10 65 14
rect 49 9 69 10
rect 49 6 69 7
rect 53 2 69 6
<< ndcontact >>
rect 22 1008 26 1012
rect 22 1000 26 1004
rect 21 980 25 984
rect 27 972 31 976
rect 27 963 31 967
rect 856 938 906 942
rect 856 930 906 934
rect 856 922 906 926
rect 57 918 77 922
rect 856 914 906 918
rect 57 910 77 914
rect 856 906 906 910
rect 57 902 77 906
rect 856 898 906 902
rect 27 874 31 878
rect 33 866 37 870
rect 849 843 889 847
rect 849 835 889 839
rect 849 827 889 831
rect 849 819 889 823
rect 849 811 889 815
rect 1151 799 1201 803
rect 22 792 26 796
rect 1151 791 1201 795
rect 22 784 26 788
rect 1633 788 1637 792
rect 1151 783 1201 787
rect 1633 780 1637 784
rect 1151 775 1201 779
rect 21 764 25 768
rect 1151 767 1201 771
rect 27 756 31 760
rect 1151 759 1201 763
rect 1632 760 1636 764
rect 27 747 31 751
rect 844 748 874 752
rect 1638 752 1642 756
rect 844 740 874 744
rect 1638 743 1642 747
rect 844 732 874 736
rect 844 724 874 728
rect 57 702 77 706
rect 57 694 77 698
rect 57 686 77 690
rect 890 674 910 678
rect 890 666 910 670
rect 27 658 31 662
rect 890 658 910 662
rect 33 650 37 654
rect 22 576 26 580
rect 851 578 891 582
rect 22 568 26 572
rect 851 570 891 574
rect 851 562 891 566
rect 21 548 25 552
rect 851 554 891 558
rect 851 546 891 550
rect 27 540 31 544
rect 27 531 31 535
rect 1157 497 1197 501
rect 846 493 876 497
rect 57 486 77 490
rect 846 485 876 489
rect 57 478 77 482
rect 1157 489 1197 493
rect 1625 488 1629 492
rect 846 477 876 481
rect 57 470 77 474
rect 1157 481 1197 485
rect 846 469 876 473
rect 1625 480 1629 484
rect 1157 473 1197 477
rect 1157 465 1197 469
rect 1624 460 1628 464
rect 1630 452 1634 456
rect 27 442 31 446
rect 1630 443 1634 447
rect 33 434 37 438
rect 890 422 910 426
rect 890 414 910 418
rect 890 406 910 410
rect 22 360 26 364
rect 22 352 26 356
rect 1625 338 1629 342
rect 21 332 25 336
rect 847 330 877 334
rect 27 324 31 328
rect 1625 330 1629 334
rect 847 322 877 326
rect 27 315 31 319
rect 847 314 877 318
rect 1164 315 1194 319
rect 847 306 877 310
rect 1164 307 1194 311
rect 1624 310 1628 314
rect 1164 299 1194 303
rect 1630 302 1634 306
rect 1164 291 1194 295
rect 1630 293 1634 297
rect 57 270 77 274
rect 57 262 77 266
rect 57 254 77 258
rect 891 259 911 263
rect 891 251 911 255
rect 891 243 911 247
rect 27 226 31 230
rect 33 218 37 222
rect 1625 200 1629 204
rect 1625 192 1629 196
rect 889 176 909 180
rect 889 168 909 172
rect 1205 175 1225 179
rect 1624 172 1628 176
rect 889 160 909 164
rect 1205 167 1225 171
rect 1205 159 1225 163
rect 1630 164 1634 168
rect 1630 155 1634 159
rect 22 144 26 148
rect 22 136 26 140
rect 21 116 25 120
rect 27 108 31 112
rect 27 99 31 103
rect 57 54 77 58
rect 57 46 77 50
rect 57 38 77 42
rect 27 10 31 14
rect 33 2 37 6
<< pdcontact >>
rect 44 1008 48 1012
rect 60 1000 64 1004
rect 60 980 64 984
rect 46 972 50 976
rect 44 963 48 967
rect 920 938 940 942
rect 920 930 940 934
rect 23 918 43 922
rect 920 922 940 926
rect 23 910 43 914
rect 920 914 940 918
rect 23 902 43 906
rect 920 906 940 910
rect 920 898 940 902
rect 65 874 69 878
rect 49 866 53 870
rect 901 843 921 847
rect 901 835 921 839
rect 901 827 921 831
rect 901 819 921 823
rect 901 811 921 815
rect 44 792 48 796
rect 1215 799 1235 803
rect 60 784 64 788
rect 1215 791 1235 795
rect 1655 788 1659 792
rect 1215 783 1235 787
rect 1671 780 1675 784
rect 1215 775 1235 779
rect 60 764 64 768
rect 1215 767 1235 771
rect 46 756 50 760
rect 1215 759 1235 763
rect 1671 760 1675 764
rect 44 747 48 751
rect 891 748 911 752
rect 1657 752 1661 756
rect 891 740 911 744
rect 1655 743 1659 747
rect 891 732 911 736
rect 891 724 911 728
rect 23 702 43 706
rect 23 694 43 698
rect 23 686 43 690
rect 856 674 876 678
rect 856 666 876 670
rect 65 658 69 662
rect 856 658 876 662
rect 49 650 53 654
rect 44 576 48 580
rect 903 578 923 582
rect 60 568 64 572
rect 903 570 923 574
rect 903 562 923 566
rect 60 548 64 552
rect 903 554 923 558
rect 903 546 923 550
rect 46 540 50 544
rect 44 531 48 535
rect 23 486 43 490
rect 893 493 913 497
rect 1209 497 1229 501
rect 23 478 43 482
rect 893 485 913 489
rect 1209 489 1229 493
rect 1647 488 1651 492
rect 23 470 43 474
rect 893 477 913 481
rect 1209 481 1229 485
rect 1663 480 1667 484
rect 893 469 913 473
rect 1209 473 1229 477
rect 1209 465 1229 469
rect 1663 460 1667 464
rect 1649 452 1653 456
rect 65 442 69 446
rect 1647 443 1651 447
rect 49 434 53 438
rect 856 422 876 426
rect 856 414 876 418
rect 856 406 876 410
rect 44 360 48 364
rect 60 352 64 356
rect 1647 338 1651 342
rect 60 332 64 336
rect 46 324 50 328
rect 894 330 914 334
rect 1663 330 1667 334
rect 44 315 48 319
rect 894 322 914 326
rect 894 314 914 318
rect 1211 315 1231 319
rect 894 306 914 310
rect 1211 307 1231 311
rect 1663 310 1667 314
rect 1211 299 1231 303
rect 1649 302 1653 306
rect 1211 291 1231 295
rect 1647 293 1651 297
rect 23 270 43 274
rect 23 262 43 266
rect 857 259 877 263
rect 23 254 43 258
rect 857 251 877 255
rect 857 243 877 247
rect 65 226 69 230
rect 49 218 53 222
rect 1647 200 1651 204
rect 1663 192 1667 196
rect 855 176 875 180
rect 1171 175 1191 179
rect 855 168 875 172
rect 1171 167 1191 171
rect 855 160 875 164
rect 1663 172 1667 176
rect 1171 159 1191 163
rect 1649 164 1653 168
rect 1647 155 1651 159
rect 44 144 48 148
rect 60 136 64 140
rect 60 116 64 120
rect 46 108 50 112
rect 44 99 48 103
rect 23 54 43 58
rect 23 46 43 50
rect 23 38 43 42
rect 65 10 69 14
rect 49 2 53 6
<< polysilicon >>
rect 18 1005 22 1007
rect 32 1005 44 1007
rect 64 1005 68 1007
rect 18 977 21 979
rect 31 977 44 979
rect 64 977 67 979
rect 14 969 15 970
rect 19 969 21 970
rect 14 968 21 969
rect 31 968 35 970
rect 38 968 44 970
rect 64 968 76 970
rect 848 935 856 937
rect 906 935 920 937
rect 940 935 943 937
rect 848 927 856 929
rect 906 927 920 929
rect 940 927 943 929
rect 848 919 856 921
rect 906 919 920 921
rect 940 919 943 921
rect 10 915 23 917
rect 43 915 57 917
rect 77 915 82 917
rect 848 911 856 913
rect 906 911 920 913
rect 940 911 943 913
rect 10 907 23 909
rect 43 907 57 909
rect 77 907 82 909
rect 848 903 856 905
rect 906 903 920 905
rect 940 903 943 905
rect 23 871 27 873
rect 37 871 49 873
rect 69 871 73 873
rect 844 840 849 842
rect 889 840 901 842
rect 921 840 924 842
rect 844 832 849 834
rect 889 832 901 834
rect 921 832 924 834
rect 844 824 849 826
rect 889 824 901 826
rect 921 824 924 826
rect 844 816 849 818
rect 889 816 901 818
rect 921 816 924 818
rect 1143 796 1151 798
rect 1201 796 1215 798
rect 1235 796 1238 798
rect 18 789 22 791
rect 32 789 44 791
rect 64 789 68 791
rect 1143 788 1151 790
rect 1201 788 1215 790
rect 1235 788 1238 790
rect 1629 785 1633 787
rect 1643 785 1655 787
rect 1675 785 1679 787
rect 1143 780 1151 782
rect 1201 780 1215 782
rect 1235 780 1238 782
rect 1143 772 1151 774
rect 1201 772 1215 774
rect 1235 772 1238 774
rect 1143 764 1151 766
rect 1201 764 1215 766
rect 1235 764 1238 766
rect 18 761 21 763
rect 31 761 44 763
rect 64 761 67 763
rect 14 753 15 754
rect 1629 757 1632 759
rect 1642 757 1655 759
rect 1675 757 1678 759
rect 19 753 21 754
rect 14 752 21 753
rect 31 752 35 754
rect 38 752 44 754
rect 64 752 76 754
rect 1625 749 1626 750
rect 1630 749 1632 750
rect 1625 748 1632 749
rect 1642 748 1646 750
rect 1649 748 1655 750
rect 1675 748 1687 750
rect 841 745 844 747
rect 874 745 891 747
rect 911 745 914 747
rect 841 737 844 739
rect 874 737 891 739
rect 911 737 914 739
rect 841 729 844 731
rect 874 729 891 731
rect 911 729 914 731
rect 10 699 23 701
rect 43 699 57 701
rect 77 699 82 701
rect 10 691 23 693
rect 43 691 57 693
rect 77 691 82 693
rect 843 671 856 673
rect 876 671 890 673
rect 910 671 915 673
rect 843 663 856 665
rect 876 663 890 665
rect 910 663 915 665
rect 23 655 27 657
rect 37 655 49 657
rect 69 655 73 657
rect 18 573 22 575
rect 32 573 44 575
rect 64 573 68 575
rect 846 575 851 577
rect 891 575 903 577
rect 923 575 926 577
rect 846 567 851 569
rect 891 567 903 569
rect 923 567 926 569
rect 846 559 851 561
rect 891 559 903 561
rect 923 559 926 561
rect 846 551 851 553
rect 891 551 903 553
rect 923 551 926 553
rect 18 545 21 547
rect 31 545 44 547
rect 64 545 67 547
rect 14 537 15 538
rect 19 537 21 538
rect 14 536 21 537
rect 31 536 35 538
rect 38 536 44 538
rect 64 536 76 538
rect 1152 494 1157 496
rect 1197 494 1209 496
rect 1229 494 1232 496
rect 843 490 846 492
rect 876 490 893 492
rect 913 490 916 492
rect 10 483 23 485
rect 43 483 57 485
rect 77 483 82 485
rect 1152 486 1157 488
rect 1197 486 1209 488
rect 1229 486 1232 488
rect 843 482 846 484
rect 876 482 893 484
rect 913 482 916 484
rect 10 475 23 477
rect 43 475 57 477
rect 77 475 82 477
rect 843 474 846 476
rect 876 474 893 476
rect 913 474 916 476
rect 1621 485 1625 487
rect 1635 485 1647 487
rect 1667 485 1671 487
rect 1152 478 1157 480
rect 1197 478 1209 480
rect 1229 478 1232 480
rect 1152 470 1157 472
rect 1197 470 1209 472
rect 1229 470 1232 472
rect 1621 457 1624 459
rect 1634 457 1647 459
rect 1667 457 1670 459
rect 1617 449 1618 450
rect 1622 449 1624 450
rect 1617 448 1624 449
rect 1634 448 1638 450
rect 1641 448 1647 450
rect 1667 448 1679 450
rect 23 439 27 441
rect 37 439 49 441
rect 69 439 73 441
rect 843 419 856 421
rect 876 419 890 421
rect 910 419 915 421
rect 843 411 856 413
rect 876 411 890 413
rect 910 411 915 413
rect 18 357 22 359
rect 32 357 44 359
rect 64 357 68 359
rect 1621 335 1625 337
rect 1635 335 1647 337
rect 1667 335 1671 337
rect 18 329 21 331
rect 31 329 44 331
rect 64 329 67 331
rect 14 321 15 322
rect 844 327 847 329
rect 877 327 894 329
rect 914 327 917 329
rect 19 321 21 322
rect 14 320 21 321
rect 31 320 35 322
rect 38 320 44 322
rect 64 320 76 322
rect 844 319 847 321
rect 877 319 894 321
rect 914 319 917 321
rect 844 311 847 313
rect 877 311 894 313
rect 914 311 917 313
rect 1161 312 1164 314
rect 1194 312 1211 314
rect 1231 312 1234 314
rect 1621 307 1624 309
rect 1634 307 1647 309
rect 1667 307 1670 309
rect 1161 304 1164 306
rect 1194 304 1211 306
rect 1231 304 1234 306
rect 1617 299 1618 300
rect 1622 299 1624 300
rect 1617 298 1624 299
rect 1634 298 1638 300
rect 1641 298 1647 300
rect 1667 298 1679 300
rect 1161 296 1164 298
rect 1194 296 1211 298
rect 1231 296 1234 298
rect 10 267 23 269
rect 43 267 57 269
rect 77 267 82 269
rect 10 259 23 261
rect 43 259 57 261
rect 77 259 82 261
rect 844 256 857 258
rect 877 256 891 258
rect 911 256 916 258
rect 844 248 857 250
rect 877 248 891 250
rect 911 248 916 250
rect 23 223 27 225
rect 37 223 49 225
rect 69 223 73 225
rect 1621 197 1625 199
rect 1635 197 1647 199
rect 1667 197 1671 199
rect 842 173 855 175
rect 875 173 889 175
rect 909 173 914 175
rect 1158 172 1171 174
rect 1191 172 1205 174
rect 1225 172 1230 174
rect 842 165 855 167
rect 875 165 889 167
rect 909 165 914 167
rect 1621 169 1624 171
rect 1634 169 1647 171
rect 1667 169 1670 171
rect 1158 164 1171 166
rect 1191 164 1205 166
rect 1225 164 1230 166
rect 1617 161 1618 162
rect 1622 161 1624 162
rect 1617 160 1624 161
rect 1634 160 1638 162
rect 1641 160 1647 162
rect 1667 160 1679 162
rect 18 141 22 143
rect 32 141 44 143
rect 64 141 68 143
rect 18 113 21 115
rect 31 113 44 115
rect 64 113 67 115
rect 14 105 15 106
rect 19 105 21 106
rect 14 104 21 105
rect 31 104 35 106
rect 38 104 44 106
rect 64 104 76 106
rect 10 51 23 53
rect 43 51 57 53
rect 77 51 82 53
rect 10 43 23 45
rect 43 43 57 45
rect 77 43 82 45
rect 23 7 27 9
rect 37 7 49 9
rect 69 7 73 9
<< polycontact >>
rect 33 1001 37 1005
rect 33 979 37 983
rect 15 969 19 973
rect 71 970 75 974
rect 844 934 848 938
rect 844 926 848 930
rect 6 914 10 918
rect 844 918 848 922
rect 6 906 10 910
rect 844 910 848 914
rect 844 902 848 906
rect 38 873 42 877
rect 840 839 844 843
rect 840 831 844 835
rect 840 823 844 827
rect 840 815 844 819
rect 1139 795 1143 799
rect 33 785 37 789
rect 1139 787 1143 791
rect 1139 779 1143 783
rect 1644 781 1648 785
rect 1139 771 1143 775
rect 33 763 37 767
rect 1139 763 1143 767
rect 15 753 19 757
rect 1644 759 1648 763
rect 71 754 75 758
rect 837 744 841 748
rect 1626 749 1630 753
rect 1682 750 1686 754
rect 837 736 841 740
rect 837 728 841 732
rect 6 698 10 702
rect 6 690 10 694
rect 839 670 843 674
rect 839 662 843 666
rect 38 657 42 661
rect 842 574 846 578
rect 33 569 37 573
rect 842 566 846 570
rect 842 558 846 562
rect 33 547 37 551
rect 842 550 846 554
rect 15 537 19 541
rect 71 538 75 542
rect 6 482 10 486
rect 839 489 843 493
rect 1148 493 1152 497
rect 6 474 10 478
rect 839 481 843 485
rect 1148 485 1152 489
rect 839 473 843 477
rect 1148 477 1152 481
rect 1636 481 1640 485
rect 1148 469 1152 473
rect 1636 459 1640 463
rect 1618 449 1622 453
rect 1674 450 1678 454
rect 38 441 42 445
rect 839 418 843 422
rect 839 410 843 414
rect 33 353 37 357
rect 33 331 37 335
rect 15 321 19 325
rect 840 326 844 330
rect 1636 331 1640 335
rect 71 322 75 326
rect 840 318 844 322
rect 840 310 844 314
rect 1157 311 1161 315
rect 1157 303 1161 307
rect 1636 309 1640 313
rect 1157 295 1161 299
rect 1618 299 1622 303
rect 1674 300 1678 304
rect 6 266 10 270
rect 6 258 10 262
rect 840 255 844 259
rect 840 247 844 251
rect 38 225 42 229
rect 1636 193 1640 197
rect 838 172 842 176
rect 838 164 842 168
rect 1154 171 1158 175
rect 1154 163 1158 167
rect 1636 171 1640 175
rect 1618 161 1622 165
rect 1674 162 1678 166
rect 33 137 37 141
rect 33 115 37 119
rect 15 105 19 109
rect 71 106 75 110
rect 6 50 10 54
rect 6 42 10 46
rect 38 9 42 13
<< metal1 >>
rect 208 1084 1498 1089
rect 192 1076 1481 1081
rect 178 1064 1466 1069
rect 155 1056 158 1061
rect 163 1056 1450 1061
rect 146 1048 1433 1053
rect 14 1010 17 1019
rect 73 1018 76 1019
rect 23 1012 28 1013
rect 73 1013 108 1018
rect -4 1007 17 1010
rect 26 1009 44 1012
rect 14 1004 17 1007
rect 73 1005 76 1013
rect 103 1010 108 1013
rect 103 1005 1697 1010
rect 34 997 37 1001
rect 64 1000 71 1004
rect -4 994 64 997
rect -4 993 -1 994
rect -13 990 -1 993
rect -44 928 -23 931
rect -44 915 -20 919
rect -24 910 -20 915
rect -13 910 -10 990
rect 20 985 24 990
rect 61 989 64 994
rect 968 993 973 1005
rect 61 986 74 989
rect 15 984 24 985
rect -3 981 11 984
rect -3 933 0 981
rect 8 959 11 981
rect 15 973 18 984
rect 33 983 36 986
rect 61 984 64 986
rect 31 972 38 975
rect 43 972 46 975
rect 71 974 74 986
rect 84 985 206 988
rect 31 964 44 967
rect 34 960 37 964
rect 907 965 1072 970
rect 8 956 15 959
rect 12 952 15 956
rect 35 955 37 960
rect 34 952 37 955
rect 909 957 913 965
rect 12 949 37 952
rect 39 937 81 940
rect -3 918 0 928
rect 14 922 18 928
rect 14 918 23 922
rect 77 918 81 937
rect 209 939 571 940
rect 209 936 844 939
rect 906 938 908 942
rect 940 938 942 942
rect 567 934 844 936
rect -3 915 6 918
rect 2 914 6 915
rect -24 906 6 910
rect 14 906 18 918
rect 93 915 296 918
rect 43 910 53 914
rect 49 906 53 910
rect 14 897 23 906
rect 49 902 57 906
rect 17 895 23 897
rect 19 893 31 895
rect 20 892 31 893
rect 49 892 53 902
rect 13 885 16 887
rect 39 888 53 892
rect 13 882 22 885
rect 19 878 22 882
rect 19 875 27 878
rect 19 862 22 875
rect 39 877 42 888
rect 77 883 79 888
rect 76 878 79 883
rect 69 875 79 878
rect 37 866 49 869
rect 39 855 42 866
rect 76 865 79 875
rect 76 859 79 860
rect 93 855 96 915
rect 39 852 96 855
rect 567 843 571 934
rect 591 926 844 931
rect 919 930 920 934
rect 612 918 844 923
rect 940 922 942 926
rect 657 913 844 914
rect 630 909 844 913
rect 919 914 920 918
rect 630 905 695 909
rect 940 906 942 910
rect 830 901 844 906
rect 851 898 856 902
rect 851 887 855 898
rect 919 898 920 902
rect 851 883 991 887
rect 892 857 1053 862
rect 892 847 896 857
rect 889 843 896 847
rect 921 843 968 847
rect 567 839 840 843
rect 892 839 896 843
rect 14 794 17 803
rect 23 796 28 797
rect 73 801 76 803
rect 73 798 84 801
rect -4 791 17 794
rect 26 793 44 796
rect 14 788 17 791
rect 73 789 76 798
rect 34 781 37 785
rect 64 784 71 788
rect -4 778 64 781
rect -4 777 -1 778
rect -13 774 -1 777
rect -42 712 -23 715
rect -42 699 -20 703
rect -24 694 -20 699
rect -13 694 -10 774
rect 20 769 24 774
rect 61 773 64 778
rect 61 770 74 773
rect 15 768 24 769
rect -3 765 11 768
rect -3 717 0 765
rect 8 743 11 765
rect 15 757 18 768
rect 33 767 36 770
rect 61 768 64 770
rect 31 756 38 759
rect 43 756 46 759
rect 71 758 74 770
rect 84 769 189 772
rect 31 748 44 751
rect 34 744 37 748
rect 567 747 571 839
rect 892 835 901 839
rect 837 834 840 835
rect 612 831 840 834
rect 837 826 840 827
rect 630 823 840 826
rect 892 823 896 835
rect 927 831 931 843
rect 921 827 931 831
rect 892 819 901 823
rect 830 816 840 819
rect 837 815 840 816
rect 927 815 931 827
rect 847 811 849 815
rect 921 811 931 815
rect 847 803 850 811
rect 847 800 992 803
rect 1048 792 1053 857
rect 1067 800 1072 965
rect 1388 850 1643 857
rect 1067 795 1139 800
rect 1201 799 1203 803
rect 1235 799 1237 803
rect 1048 787 1139 792
rect 1214 791 1215 795
rect 1006 780 1139 784
rect 1235 783 1237 787
rect 885 779 1139 780
rect 885 777 1012 779
rect 1040 770 1139 775
rect 1214 775 1215 779
rect 874 748 880 752
rect 911 748 920 752
rect 1040 750 1045 770
rect 1235 767 1237 771
rect 8 740 15 743
rect 12 736 15 740
rect 35 739 37 744
rect 34 736 37 739
rect 12 733 37 736
rect 567 744 837 747
rect 880 744 884 748
rect 39 721 81 724
rect -3 702 0 712
rect 14 706 18 712
rect 14 702 23 706
rect 77 702 81 721
rect -3 699 6 702
rect 2 698 6 699
rect -24 690 6 694
rect 14 690 18 702
rect 93 699 278 702
rect 43 694 53 698
rect 49 690 53 694
rect 14 681 23 690
rect 49 686 57 690
rect 17 679 23 681
rect 19 677 31 679
rect 20 676 31 677
rect 49 676 53 686
rect 13 669 16 671
rect 39 672 53 676
rect 13 666 22 669
rect 19 662 22 666
rect 19 659 27 662
rect 19 643 22 659
rect 39 661 42 672
rect 77 667 79 672
rect 76 662 79 667
rect 69 659 79 662
rect 37 650 49 653
rect 39 639 42 650
rect 76 649 79 659
rect 76 643 79 644
rect 93 639 96 699
rect 567 674 571 744
rect 880 740 891 744
rect 613 736 837 739
rect 691 728 837 731
rect 882 728 886 740
rect 916 736 920 748
rect 911 732 920 736
rect 916 730 920 732
rect 882 724 891 728
rect 916 726 969 730
rect 855 714 859 724
rect 855 710 990 714
rect 847 686 969 690
rect 847 678 851 686
rect 910 679 990 683
rect 847 674 856 678
rect 910 674 914 679
rect 567 670 839 674
rect 648 663 656 664
rect 663 663 839 666
rect 648 662 839 663
rect 847 662 851 674
rect 876 666 886 670
rect 882 662 886 666
rect 648 659 667 662
rect 648 656 656 659
rect 847 658 856 662
rect 882 658 890 662
rect 882 654 886 658
rect 1041 654 1045 750
rect 882 650 1045 654
rect 1058 762 1139 767
rect 1388 773 1395 850
rect 1692 799 1697 1005
rect 1742 850 1759 857
rect 1625 783 1628 799
rect 1634 792 1639 793
rect 1684 796 1700 799
rect 1637 789 1655 792
rect 1614 780 1633 783
rect 1684 784 1687 796
rect 1692 795 1700 796
rect 1645 777 1648 781
rect 1675 780 1687 784
rect 1502 774 1675 777
rect 1302 769 1395 773
rect 1388 768 1395 769
rect 1631 765 1635 770
rect 1672 769 1675 774
rect 1672 766 1685 769
rect 1626 764 1635 765
rect 1058 646 1063 762
rect 1146 759 1151 763
rect 1146 751 1150 759
rect 1214 759 1215 763
rect 1626 753 1629 764
rect 1644 763 1647 766
rect 1672 764 1675 766
rect 1642 752 1649 755
rect 1654 752 1657 755
rect 1682 754 1685 766
rect 1642 744 1655 747
rect 1645 740 1648 744
rect 39 636 96 639
rect 301 638 1063 646
rect 1391 735 1641 739
rect 1646 735 1648 740
rect 894 592 1112 596
rect 14 578 17 587
rect 73 586 76 587
rect 23 580 28 581
rect 73 583 83 586
rect -4 575 17 578
rect 26 577 44 580
rect 14 572 17 575
rect 73 573 76 583
rect 894 582 898 592
rect 891 578 898 582
rect 923 578 969 582
rect 664 575 842 578
rect 34 565 37 569
rect 64 568 71 572
rect 193 574 842 575
rect 894 574 898 578
rect 193 569 554 574
rect 559 570 675 574
rect 894 570 903 574
rect 559 569 655 570
rect 664 569 675 570
rect -4 562 64 565
rect -4 561 -1 562
rect -13 558 -1 561
rect -42 496 -23 499
rect -42 483 -20 487
rect -24 478 -20 483
rect -13 478 -10 558
rect 20 553 24 558
rect 61 557 64 562
rect 611 558 662 561
rect 61 554 74 557
rect 15 552 24 553
rect -3 549 11 552
rect -3 501 0 549
rect 8 527 11 549
rect 15 541 18 552
rect 33 551 36 554
rect 61 552 64 554
rect 31 540 38 543
rect 43 540 46 543
rect 71 542 74 554
rect 84 553 174 556
rect 659 549 663 550
rect 627 546 663 549
rect 31 532 44 535
rect 34 528 37 532
rect 8 524 15 527
rect 12 520 15 524
rect 35 523 37 528
rect 34 520 37 523
rect 12 517 37 520
rect 39 505 81 508
rect -3 486 0 496
rect 14 490 18 496
rect 14 486 23 490
rect 77 486 81 505
rect 669 492 675 569
rect 699 567 842 570
rect 699 564 702 567
rect 839 566 842 567
rect 683 561 702 564
rect 709 559 842 562
rect 709 553 712 559
rect 839 558 842 559
rect 894 558 898 570
rect 929 566 933 578
rect 923 562 933 566
rect 683 550 712 553
rect 894 554 903 558
rect 825 551 842 554
rect 839 550 842 551
rect 929 550 933 562
rect 849 546 851 550
rect 923 546 933 550
rect 849 535 852 546
rect 849 532 991 535
rect 947 505 1055 508
rect 876 493 882 497
rect 913 493 922 497
rect 669 489 839 492
rect 882 489 886 493
rect -3 483 6 486
rect 2 482 6 483
rect -24 474 6 478
rect 14 474 18 486
rect 93 483 263 486
rect 611 483 659 486
rect 43 478 53 482
rect 49 474 53 478
rect 14 465 23 474
rect 49 470 57 474
rect 17 463 23 465
rect 19 461 31 463
rect 20 460 31 461
rect 49 460 53 470
rect 13 453 16 455
rect 39 456 53 460
rect 13 450 22 453
rect 19 446 22 450
rect 19 443 27 446
rect 19 427 22 443
rect 39 445 42 456
rect 77 451 79 456
rect 76 446 79 451
rect 69 443 79 446
rect 37 434 49 437
rect 39 423 42 434
rect 76 433 79 443
rect 76 427 79 428
rect 93 423 96 483
rect 39 420 96 423
rect 669 422 675 489
rect 882 485 893 489
rect 683 481 839 484
rect 835 473 839 476
rect 884 473 888 485
rect 918 481 922 493
rect 1052 488 1055 505
rect 1108 497 1112 592
rect 1200 515 1275 519
rect 1200 501 1204 515
rect 1197 497 1204 501
rect 1229 497 1247 501
rect 1108 493 1148 497
rect 1200 493 1204 497
rect 1200 489 1209 493
rect 1145 488 1148 489
rect 1052 485 1148 488
rect 913 477 922 481
rect 1145 480 1148 481
rect 918 473 967 477
rect 1021 477 1148 480
rect 1200 477 1204 489
rect 1235 485 1239 497
rect 1229 481 1239 485
rect 884 469 893 473
rect 918 471 922 473
rect 857 462 861 469
rect 857 458 990 462
rect 847 434 969 438
rect 847 426 851 434
rect 910 430 914 431
rect 910 426 990 430
rect 847 422 856 426
rect 910 422 914 426
rect 669 418 839 422
rect 693 407 832 411
rect 835 407 839 414
rect 847 410 851 422
rect 876 414 886 418
rect 882 410 886 414
rect 693 403 839 407
rect 847 406 856 410
rect 882 406 890 410
rect 882 396 886 406
rect 1021 396 1024 477
rect 1200 473 1209 477
rect 1145 472 1148 473
rect 1112 469 1148 472
rect 1235 469 1239 481
rect 882 392 1027 396
rect 1112 385 1115 469
rect 1155 465 1157 469
rect 1229 465 1239 469
rect 1155 461 1158 465
rect 1243 446 1247 497
rect 1271 476 1275 515
rect 1391 476 1395 735
rect 1615 726 1625 731
rect 1622 509 1625 726
rect 1697 524 1700 795
rect 1716 769 1725 772
rect 1617 506 1625 509
rect 1689 521 1700 524
rect 1617 483 1620 506
rect 1689 499 1692 521
rect 1626 492 1631 493
rect 1676 496 1692 499
rect 1629 489 1647 492
rect 1606 480 1625 483
rect 1676 484 1679 496
rect 1271 472 1395 476
rect 1637 477 1640 481
rect 1667 480 1679 484
rect 1485 474 1667 477
rect 1623 465 1627 470
rect 1664 469 1667 474
rect 1664 466 1677 469
rect 1618 464 1627 465
rect 1618 453 1621 464
rect 1636 463 1639 466
rect 1664 464 1667 466
rect 1634 452 1641 455
rect 1646 452 1649 455
rect 1674 454 1677 466
rect 1634 444 1647 447
rect 1637 440 1640 444
rect 1391 435 1633 439
rect 1638 435 1640 440
rect 284 377 640 385
rect 648 377 1119 385
rect 14 362 17 371
rect 23 364 28 365
rect 73 369 76 371
rect 73 366 84 369
rect -4 359 17 362
rect 26 361 44 364
rect 14 356 17 359
rect 73 357 76 366
rect 34 349 37 353
rect 64 352 71 356
rect -4 346 64 349
rect -4 345 -1 346
rect -13 342 -1 345
rect -39 280 -23 283
rect -39 267 -20 271
rect -24 262 -20 267
rect -13 262 -10 342
rect 20 337 24 342
rect 61 341 64 346
rect 946 344 1124 347
rect 61 338 74 341
rect 15 336 24 337
rect -3 333 11 336
rect -3 285 0 333
rect 8 311 11 333
rect 15 325 18 336
rect 33 335 36 338
rect 61 336 64 338
rect 31 324 38 327
rect 43 324 46 327
rect 71 326 74 338
rect 84 337 157 340
rect 877 330 883 334
rect 914 330 923 334
rect 176 324 607 329
rect 612 326 840 329
rect 883 326 887 330
rect 612 324 781 326
rect 31 316 44 319
rect 34 312 37 316
rect 8 308 15 311
rect 12 304 15 308
rect 35 307 37 312
rect 34 304 37 307
rect 12 301 37 304
rect 39 289 81 292
rect -3 270 0 280
rect 14 274 18 280
rect 14 270 23 274
rect 77 270 81 289
rect -3 267 6 270
rect 2 266 6 267
rect -24 258 6 262
rect 14 258 18 270
rect 93 267 248 270
rect 43 262 53 266
rect 49 258 53 262
rect 14 249 23 258
rect 49 254 57 258
rect 17 247 23 249
rect 19 245 31 247
rect 20 244 31 245
rect 49 244 53 254
rect 13 237 16 239
rect 39 240 53 244
rect 13 234 22 237
rect 19 230 22 234
rect 19 227 27 230
rect 19 211 22 227
rect 39 229 42 240
rect 77 235 79 240
rect 76 230 79 235
rect 69 227 79 230
rect 37 218 49 221
rect 39 207 42 218
rect 76 217 79 227
rect 76 211 79 212
rect 93 207 96 267
rect 703 259 707 324
rect 883 322 894 326
rect 713 318 840 321
rect 713 299 716 318
rect 825 310 840 313
rect 885 310 889 322
rect 919 318 923 330
rect 914 314 923 318
rect 919 312 923 314
rect 1120 314 1124 344
rect 1194 315 1200 319
rect 1231 315 1240 319
rect 885 306 894 310
rect 919 308 968 312
rect 1120 311 1157 314
rect 1200 311 1204 315
rect 1200 307 1211 311
rect 1006 306 1010 307
rect 858 297 862 306
rect 1005 303 1157 306
rect 858 293 989 297
rect 848 271 969 275
rect 848 263 852 271
rect 911 264 990 268
rect 848 259 857 263
rect 911 259 915 264
rect 703 255 840 259
rect 834 247 840 251
rect 848 247 852 259
rect 877 251 887 255
rect 883 247 887 251
rect 848 243 857 247
rect 883 243 891 247
rect 883 240 887 243
rect 1006 240 1010 303
rect 883 236 1010 240
rect 1134 295 1157 298
rect 1202 295 1206 307
rect 1236 303 1240 315
rect 1231 299 1240 303
rect 1391 304 1395 435
rect 1607 426 1617 431
rect 1614 366 1617 426
rect 1614 358 1620 366
rect 1617 333 1620 358
rect 1689 349 1692 496
rect 1708 469 1717 472
rect 1626 342 1631 343
rect 1676 346 1692 349
rect 1629 339 1647 342
rect 1606 330 1625 333
rect 1676 334 1679 346
rect 1637 327 1640 331
rect 1667 330 1679 334
rect 1472 324 1667 327
rect 1268 301 1395 304
rect 1623 315 1627 320
rect 1664 319 1667 324
rect 1664 316 1677 319
rect 1618 314 1627 315
rect 1618 303 1621 314
rect 1636 313 1639 316
rect 1664 314 1667 316
rect 1634 302 1641 305
rect 1646 302 1649 305
rect 1674 304 1677 316
rect 1134 228 1137 295
rect 1202 291 1211 295
rect 1175 286 1179 291
rect 1236 276 1240 299
rect 1634 294 1647 297
rect 1637 290 1640 294
rect 1383 285 1633 289
rect 1638 285 1640 290
rect 269 220 685 228
rect 693 220 1141 228
rect 1134 219 1137 220
rect 39 204 96 207
rect 846 189 969 193
rect 995 192 1025 196
rect 846 180 850 189
rect 1021 188 1229 192
rect 909 184 913 185
rect 909 180 991 184
rect 1056 181 1166 185
rect 846 176 855 180
rect 909 176 913 180
rect 163 165 622 173
rect 630 171 680 173
rect 685 172 838 176
rect 685 171 689 172
rect 630 167 689 171
rect 630 165 680 167
rect 818 164 838 168
rect 846 164 850 176
rect 1056 176 1060 181
rect 1162 179 1166 181
rect 973 172 1060 176
rect 1107 173 1154 177
rect 1162 175 1171 179
rect 1225 175 1229 188
rect 875 168 885 172
rect 881 164 885 168
rect 14 146 17 155
rect 23 148 28 149
rect 73 152 76 155
rect 73 149 84 152
rect -4 143 17 146
rect 26 145 44 148
rect 14 140 17 143
rect 73 141 76 149
rect 34 133 37 137
rect 64 136 71 140
rect 818 133 822 164
rect 846 160 855 164
rect 881 160 889 164
rect 881 153 885 160
rect 1107 153 1111 173
rect 1150 171 1154 173
rect 881 149 1111 153
rect 1134 163 1154 167
rect 1162 163 1166 175
rect 1383 171 1387 285
rect 1607 276 1617 281
rect 1614 225 1617 276
rect 1614 222 1620 225
rect 1617 195 1620 222
rect 1689 211 1692 346
rect 1708 319 1717 322
rect 1626 204 1631 205
rect 1676 208 1692 211
rect 1629 201 1647 204
rect 1606 192 1625 195
rect 1676 196 1679 208
rect 1637 189 1640 193
rect 1667 192 1679 196
rect 1453 186 1667 189
rect 1191 167 1201 171
rect 1239 168 1387 171
rect 1623 177 1627 182
rect 1664 181 1667 186
rect 1664 178 1677 181
rect 1618 176 1627 177
rect 1239 167 1386 168
rect 1197 163 1201 167
rect 1134 133 1138 163
rect 1162 159 1171 163
rect 1197 159 1205 163
rect 1197 153 1201 159
rect 1239 153 1243 167
rect 1618 165 1621 176
rect 1636 175 1639 178
rect 1664 176 1667 178
rect 1634 164 1641 167
rect 1646 164 1649 167
rect 1674 166 1677 178
rect 1634 156 1647 159
rect 1197 149 1243 153
rect 1637 152 1640 156
rect 1379 147 1633 151
rect 1638 147 1640 152
rect -4 130 64 133
rect -4 129 -1 130
rect -13 126 -1 129
rect -40 64 -23 67
rect -40 51 -20 55
rect -24 46 -20 51
rect -13 46 -10 126
rect 20 121 24 126
rect 61 125 64 130
rect 61 122 74 125
rect 15 120 24 121
rect -3 117 11 120
rect -3 69 0 117
rect 8 95 11 117
rect 15 109 18 120
rect 33 119 36 122
rect 61 120 64 122
rect 31 108 38 111
rect 43 108 46 111
rect 71 110 74 122
rect 84 121 141 124
rect 254 132 1139 133
rect 254 127 678 132
rect 683 127 1139 132
rect 254 125 1139 127
rect 31 100 44 103
rect 34 96 37 100
rect 8 92 15 95
rect 12 88 15 92
rect 35 91 37 96
rect 34 88 37 91
rect 12 85 37 88
rect 237 91 680 93
rect 818 91 822 125
rect 1379 91 1383 147
rect 1607 138 1617 143
rect 237 87 1387 91
rect 237 85 680 87
rect 729 86 733 87
rect 1440 79 1573 86
rect 39 73 106 76
rect 77 72 106 73
rect -3 54 0 64
rect 14 58 18 64
rect 14 54 23 58
rect 77 54 81 72
rect -3 51 6 54
rect 2 50 6 51
rect -24 42 6 46
rect 14 42 18 54
rect 93 51 232 54
rect 1614 54 1617 138
rect 1689 126 1692 208
rect 1708 181 1717 184
rect 1665 79 1718 86
rect 1398 51 1617 54
rect 43 46 53 50
rect 49 42 53 46
rect 14 33 23 42
rect 49 38 57 42
rect 17 31 23 33
rect 19 29 31 31
rect 20 28 31 29
rect 49 28 53 38
rect 13 21 16 23
rect 39 24 53 28
rect 13 18 22 21
rect 19 14 22 18
rect 19 11 27 14
rect 19 -5 22 11
rect 39 13 42 24
rect 77 19 79 24
rect 76 14 79 19
rect 69 11 79 14
rect 37 2 49 5
rect 39 -9 42 2
rect 76 1 79 11
rect 76 -5 79 -4
rect 93 -9 96 51
rect 989 -6 995 12
rect 114 -7 1076 -6
rect 1398 -7 1401 51
rect 39 -12 96 -9
rect 114 -9 1401 -7
rect 111 -10 1401 -9
rect 111 -12 1076 -10
rect 111 -13 118 -12
<< m2contact >>
rect 203 1084 208 1089
rect 1498 1084 1503 1089
rect 187 1076 192 1081
rect 1481 1076 1486 1081
rect 173 1064 178 1069
rect 1466 1064 1471 1069
rect 158 1056 163 1061
rect 1450 1056 1455 1061
rect 141 1048 146 1053
rect 1433 1048 1438 1053
rect 23 1013 28 1018
rect -9 1005 -4 1010
rect 71 1000 76 1005
rect -23 927 -18 932
rect 15 985 20 990
rect 38 971 43 976
rect 79 984 84 989
rect 206 985 211 990
rect 968 988 973 993
rect 909 952 914 957
rect 34 936 39 941
rect -3 928 2 933
rect 204 936 209 941
rect 908 938 913 943
rect 942 937 947 942
rect 296 915 301 920
rect 11 887 16 892
rect 31 891 36 896
rect 72 883 77 888
rect 19 857 24 862
rect 75 860 80 865
rect 586 926 591 931
rect 914 929 919 934
rect 607 918 612 923
rect 942 921 947 926
rect 622 905 630 913
rect 914 913 919 918
rect 825 901 830 906
rect 942 905 947 910
rect 914 897 919 902
rect 991 883 996 888
rect 968 843 973 848
rect 23 797 28 802
rect -9 789 -4 794
rect 84 797 89 802
rect 71 784 76 789
rect -23 711 -18 716
rect 15 769 20 774
rect 38 755 43 760
rect 79 768 84 773
rect 189 769 194 774
rect 607 831 612 836
rect 625 823 630 828
rect 825 815 830 820
rect 992 800 997 805
rect 1643 850 1650 857
rect 1203 799 1208 804
rect 1237 798 1242 803
rect 1209 790 1214 795
rect 880 776 885 781
rect 1237 782 1242 787
rect 1209 774 1214 779
rect 880 748 885 753
rect 34 720 39 725
rect -3 712 2 717
rect 278 699 283 704
rect 11 671 16 676
rect 31 675 36 680
rect 72 667 77 672
rect 75 644 80 649
rect 608 736 613 741
rect 686 728 691 733
rect 969 726 974 731
rect 990 710 995 715
rect 969 686 974 691
rect 990 679 995 684
rect 640 656 648 664
rect 1237 766 1242 771
rect 1297 769 1302 774
rect 1735 850 1742 857
rect 1609 780 1614 785
rect 1634 793 1639 798
rect 1497 773 1502 778
rect 1626 765 1631 770
rect 1209 758 1214 763
rect 1146 746 1151 751
rect 1649 751 1654 756
rect 293 638 301 646
rect 23 581 28 586
rect -9 573 -4 578
rect 83 582 88 587
rect 969 578 974 583
rect 71 568 76 573
rect 187 569 193 575
rect 554 569 559 574
rect -23 495 -18 500
rect 15 553 20 558
rect 606 558 611 563
rect 657 561 662 566
rect 38 539 43 544
rect 79 552 84 557
rect 174 553 179 558
rect 622 546 627 551
rect 34 504 39 509
rect -3 496 2 501
rect 678 560 683 565
rect 678 550 683 555
rect 820 551 825 556
rect 991 532 996 537
rect 942 504 947 509
rect 882 493 887 498
rect 263 483 268 488
rect 606 483 611 488
rect 11 455 16 460
rect 31 459 36 464
rect 72 451 77 456
rect 75 428 80 433
rect 659 482 664 487
rect 678 480 683 485
rect 830 473 835 478
rect 990 458 995 463
rect 969 434 974 439
rect 990 426 995 431
rect 685 403 693 411
rect 1155 456 1160 461
rect 1610 726 1615 731
rect 1711 768 1716 773
rect 1601 480 1606 485
rect 1626 493 1631 498
rect 1480 474 1485 479
rect 1618 465 1623 470
rect 1641 451 1646 456
rect 1243 441 1248 446
rect 276 377 284 385
rect 640 377 648 385
rect 23 365 28 370
rect -9 357 -4 362
rect 84 365 89 370
rect 71 352 76 357
rect -23 279 -18 284
rect 15 337 20 342
rect 941 343 946 348
rect 38 323 43 328
rect 79 336 84 341
rect 157 337 162 342
rect 883 330 888 335
rect 171 324 176 329
rect 607 324 612 329
rect 34 288 39 293
rect -3 280 2 285
rect 248 267 253 272
rect 11 239 16 244
rect 31 243 36 248
rect 72 235 77 240
rect 75 212 80 217
rect 820 310 825 315
rect 1200 315 1205 320
rect 968 308 973 313
rect 712 294 717 299
rect 969 271 974 276
rect 990 264 995 269
rect 829 247 834 252
rect 1263 300 1268 305
rect 1602 426 1607 431
rect 1601 330 1606 335
rect 1703 468 1708 473
rect 1626 343 1631 348
rect 1467 324 1472 329
rect 1618 315 1623 320
rect 1641 301 1646 306
rect 1175 281 1180 286
rect 1236 271 1241 276
rect 261 220 269 228
rect 685 220 693 228
rect 969 189 974 194
rect 990 192 995 197
rect 991 180 996 185
rect 155 165 163 173
rect 622 165 630 173
rect 968 172 973 177
rect 23 149 28 154
rect -9 141 -4 146
rect 84 148 89 153
rect 71 136 76 141
rect 1602 276 1607 281
rect 1601 192 1606 197
rect 1703 318 1708 323
rect 1626 205 1631 210
rect 1448 186 1453 191
rect 1618 177 1623 182
rect 1641 163 1646 168
rect -23 63 -18 68
rect 15 121 20 126
rect 38 107 43 112
rect 79 120 84 125
rect 141 121 146 126
rect 246 125 254 133
rect 678 127 683 132
rect 229 85 237 93
rect 729 91 734 96
rect 1602 138 1607 143
rect 1433 79 1440 86
rect 1573 79 1580 86
rect 34 72 39 77
rect 106 72 111 77
rect -3 64 2 69
rect 1703 180 1708 185
rect 1658 79 1665 86
rect 11 23 16 28
rect 31 27 36 32
rect 72 19 77 24
rect 75 -4 80 1
rect 989 12 995 18
rect 106 -13 111 -8
<< pdm12contact >>
rect 659 550 664 555
rect 967 473 972 478
rect 989 293 994 298
rect 232 51 237 56
<< metal2 >>
rect 140 1053 147 1093
rect 140 1048 141 1053
rect 146 1048 147 1053
rect 2 1014 23 1017
rect -14 1006 -9 1009
rect 2 990 5 1014
rect 72 999 76 1000
rect 2 987 15 990
rect 39 953 42 971
rect 79 953 82 984
rect 39 950 82 953
rect 29 938 34 941
rect -18 929 -3 932
rect 31 887 34 891
rect 31 884 72 887
rect 82 886 86 892
rect 82 883 87 886
rect -30 858 19 861
rect -30 676 -27 858
rect 84 864 87 883
rect 80 861 87 864
rect 84 802 87 861
rect 2 798 23 801
rect -14 790 -9 793
rect 2 774 5 798
rect 72 783 76 784
rect 2 771 15 774
rect 39 737 42 755
rect 79 737 82 768
rect 39 734 82 737
rect 29 722 34 725
rect -18 713 -3 716
rect 140 709 147 1048
rect 139 702 147 709
rect -30 673 11 676
rect -30 459 -27 673
rect 31 671 34 675
rect 31 668 72 671
rect 82 670 86 676
rect 82 667 87 670
rect 84 648 87 667
rect 80 645 87 648
rect 84 587 87 645
rect 2 582 23 585
rect -14 574 -9 577
rect 2 558 5 582
rect 72 567 76 568
rect 2 555 15 558
rect 39 521 42 539
rect 79 521 82 552
rect 39 518 82 521
rect 29 506 34 509
rect -18 497 -3 500
rect -34 456 11 459
rect -31 243 -28 456
rect 31 455 34 459
rect 31 452 72 455
rect 82 454 86 460
rect 82 451 87 454
rect 140 453 147 702
rect 84 432 87 451
rect 139 446 147 453
rect 80 429 87 432
rect 84 370 87 429
rect 2 366 23 369
rect -14 358 -9 361
rect 2 342 5 366
rect 72 351 76 352
rect 2 339 15 342
rect 39 305 42 323
rect 79 305 82 336
rect 39 302 82 305
rect 29 290 34 293
rect -18 281 -3 284
rect -31 240 11 243
rect -31 28 -28 240
rect 31 239 34 243
rect 31 236 72 239
rect 82 238 86 244
rect 82 235 87 238
rect 84 216 87 235
rect 80 213 87 216
rect 2 150 23 153
rect -14 142 -9 145
rect 2 126 5 150
rect 84 153 87 213
rect 140 154 147 446
rect 139 147 147 154
rect 72 135 76 136
rect 2 123 15 126
rect 140 126 147 147
rect 140 121 141 126
rect 146 121 147 126
rect 39 89 42 107
rect 79 89 82 120
rect 39 86 82 89
rect 29 74 34 77
rect -18 65 -3 68
rect -31 25 11 28
rect 31 23 34 27
rect 31 20 72 23
rect 82 22 86 28
rect 82 19 87 22
rect 84 0 87 19
rect 80 -3 87 0
rect 106 -8 110 72
rect 140 -39 147 121
rect 155 1061 162 1093
rect 172 1069 179 1094
rect 172 1064 173 1069
rect 178 1064 179 1069
rect 155 1056 158 1061
rect 155 709 162 1056
rect 172 709 179 1064
rect 187 1081 194 1095
rect 192 1076 194 1081
rect 187 774 194 1076
rect 187 769 189 774
rect 187 709 194 769
rect 203 1089 210 1094
rect 208 1084 210 1089
rect 203 990 210 1084
rect 203 985 206 990
rect 203 941 210 985
rect 203 936 204 941
rect 209 936 210 941
rect 203 709 210 936
rect 230 709 237 1095
rect 246 709 253 1095
rect 155 702 163 709
rect 171 702 179 709
rect 186 702 194 709
rect 202 702 210 709
rect 229 702 237 709
rect 245 702 253 709
rect 155 453 162 702
rect 172 558 179 702
rect 172 553 174 558
rect 172 453 179 553
rect 187 575 194 702
rect 193 569 194 575
rect 187 453 194 569
rect 203 453 210 702
rect 230 453 237 702
rect 246 453 253 702
rect 155 446 163 453
rect 171 446 179 453
rect 186 446 194 453
rect 202 446 210 453
rect 229 446 237 453
rect 245 446 253 453
rect 155 342 162 446
rect 155 337 157 342
rect 155 173 162 337
rect 172 329 179 446
rect 176 324 179 329
rect 155 154 162 165
rect 172 154 179 324
rect 187 154 194 446
rect 203 154 210 446
rect 230 154 237 446
rect 246 272 253 446
rect 246 267 248 272
rect 246 154 253 267
rect 155 147 163 154
rect 171 147 179 154
rect 186 147 194 154
rect 202 147 210 154
rect 229 147 237 154
rect 245 147 253 154
rect 155 -39 162 147
rect 172 -39 179 147
rect 187 -38 194 147
rect 203 -41 210 147
rect 230 93 237 147
rect 230 56 237 85
rect 230 51 232 56
rect 230 -41 237 51
rect 246 133 253 147
rect 261 709 268 1095
rect 276 709 283 1094
rect 293 920 300 1095
rect 1433 1053 1440 1120
rect 1438 1048 1440 1053
rect 909 943 913 952
rect 968 942 973 988
rect 909 934 913 938
rect 947 938 973 942
rect 554 926 586 931
rect 909 930 914 934
rect 293 915 296 920
rect 293 709 300 915
rect 261 702 269 709
rect 276 704 284 709
rect 261 488 268 702
rect 261 483 263 488
rect 261 453 268 483
rect 276 699 278 704
rect 283 702 284 704
rect 292 702 300 709
rect 276 453 283 699
rect 293 646 300 702
rect 293 453 300 638
rect 554 574 559 926
rect 607 836 612 918
rect 914 918 918 929
rect 942 926 946 937
rect 607 741 612 831
rect 622 828 630 905
rect 811 901 825 906
rect 914 902 918 913
rect 942 910 946 921
rect 622 823 625 828
rect 607 736 608 741
rect 607 563 612 736
rect 611 558 612 563
rect 607 488 612 558
rect 611 483 612 488
rect 261 446 269 453
rect 276 446 284 453
rect 292 446 300 453
rect 261 228 268 446
rect 276 385 283 446
rect 261 154 268 220
rect 276 154 283 377
rect 293 154 300 446
rect 607 329 612 483
rect 622 551 630 823
rect 968 848 973 938
rect 722 819 825 820
rect 721 817 825 819
rect 627 546 630 551
rect 622 305 630 546
rect 640 385 648 656
rect 662 562 678 565
rect 664 551 678 554
rect 664 482 678 485
rect 687 411 690 728
rect 721 477 725 817
rect 880 756 883 776
rect 879 753 883 756
rect 968 742 973 843
rect 989 888 995 954
rect 989 883 991 888
rect 989 805 995 883
rect 1204 818 1301 822
rect 989 800 992 805
rect 1204 804 1208 818
rect 989 750 995 800
rect 1204 795 1208 799
rect 1242 799 1251 803
rect 1204 791 1209 795
rect 1209 779 1213 790
rect 1237 787 1241 798
rect 1209 763 1213 774
rect 1237 771 1241 782
rect 989 746 1146 750
rect 968 739 983 742
rect 968 738 979 739
rect 968 731 973 738
rect 968 726 969 731
rect 968 691 973 726
rect 989 715 995 746
rect 1247 738 1251 799
rect 1297 774 1301 818
rect 1093 734 1251 738
rect 989 710 990 715
rect 968 686 969 691
rect 968 583 973 686
rect 989 684 995 710
rect 989 679 990 684
rect 968 578 969 583
rect 816 552 820 555
rect 882 504 942 507
rect 882 501 885 504
rect 881 498 885 501
rect 968 478 973 578
rect 721 474 830 477
rect 667 307 668 309
rect 685 311 693 403
rect 673 308 710 311
rect 667 305 673 307
rect 621 302 673 305
rect 622 299 673 302
rect 622 173 630 299
rect 685 228 693 308
rect 711 299 714 307
rect 711 295 712 299
rect 721 251 725 474
rect 972 473 973 478
rect 968 449 973 473
rect 989 537 995 679
rect 989 532 991 537
rect 989 463 995 532
rect 989 458 990 463
rect 995 458 1155 460
rect 989 457 1155 458
rect 968 446 982 449
rect 968 445 978 446
rect 968 439 973 445
rect 968 434 969 439
rect 883 343 941 346
rect 883 338 886 343
rect 882 335 886 338
rect 816 311 820 314
rect 968 313 973 434
rect 968 276 973 308
rect 989 431 995 457
rect 1049 441 1243 445
rect 989 426 990 431
rect 989 298 995 426
rect 1199 332 1266 335
rect 1199 323 1202 332
rect 1199 320 1203 323
rect 1263 305 1266 332
rect 994 293 995 298
rect 989 285 995 293
rect 989 281 1175 285
rect 968 271 969 276
rect 974 271 979 275
rect 706 247 829 251
rect 261 147 269 154
rect 276 147 284 154
rect 292 147 300 154
rect 246 -41 253 125
rect 261 -40 268 147
rect 276 -39 283 147
rect 293 -39 300 147
rect 706 131 710 247
rect 968 194 973 271
rect 989 269 995 281
rect 1073 271 1236 275
rect 989 264 990 269
rect 989 197 995 264
rect 968 189 969 194
rect 989 192 990 197
rect 968 177 973 189
rect 968 144 973 172
rect 989 185 995 192
rect 989 180 991 185
rect 683 127 710 131
rect 729 96 733 103
rect 989 18 995 180
rect 1433 86 1440 1048
rect 1433 -26 1440 79
rect 1448 1061 1455 1122
rect 1448 1056 1450 1061
rect 1448 191 1455 1056
rect 1453 186 1455 191
rect 1448 -26 1455 186
rect 1465 1069 1472 1123
rect 1465 1064 1466 1069
rect 1471 1064 1472 1069
rect 1465 329 1472 1064
rect 1465 324 1467 329
rect 1465 -26 1472 324
rect 1480 1081 1487 1123
rect 1480 1076 1481 1081
rect 1486 1076 1487 1081
rect 1480 479 1487 1076
rect 1485 474 1487 479
rect 1480 -26 1487 474
rect 1496 1089 1503 1122
rect 1496 1084 1498 1089
rect 1496 778 1503 1084
rect 1650 850 1735 857
rect 1621 794 1634 797
rect 1496 773 1497 778
rect 1502 773 1503 778
rect 1496 -26 1503 773
rect 1610 731 1613 780
rect 1621 770 1624 794
rect 1621 767 1626 770
rect 1691 768 1711 771
rect 1650 735 1653 751
rect 1691 735 1694 768
rect 1650 732 1694 735
rect 1613 494 1626 497
rect 1602 431 1605 480
rect 1613 470 1616 494
rect 1613 467 1618 470
rect 1683 468 1703 471
rect 1642 435 1645 451
rect 1683 435 1686 468
rect 1642 432 1686 435
rect 1613 344 1626 347
rect 1602 281 1605 330
rect 1613 320 1616 344
rect 1613 317 1618 320
rect 1683 318 1703 321
rect 1642 285 1645 301
rect 1683 285 1686 318
rect 1642 282 1686 285
rect 1613 206 1626 209
rect 1602 143 1605 192
rect 1613 182 1616 206
rect 1613 179 1618 182
rect 1683 180 1703 183
rect 1642 147 1645 163
rect 1683 147 1686 180
rect 1642 144 1686 147
rect 1580 79 1658 86
<< m3contact >>
rect -19 1005 -14 1010
rect 72 994 77 999
rect 24 937 29 942
rect 16 887 21 892
rect 82 892 87 897
rect -19 789 -14 794
rect 72 778 77 783
rect 24 721 29 726
rect 16 671 21 676
rect 82 676 87 681
rect -19 573 -14 578
rect 72 562 77 567
rect 24 505 29 510
rect 16 455 21 460
rect 82 460 87 465
rect -19 357 -14 362
rect 72 346 77 351
rect 24 289 29 294
rect 16 239 21 244
rect 82 244 87 249
rect -19 141 -14 146
rect 72 130 77 135
rect 24 73 29 78
rect 16 23 21 28
rect 82 28 87 33
rect 806 901 811 906
rect 979 734 984 739
rect 1088 734 1093 739
rect 811 551 816 556
rect 668 307 673 312
rect 710 307 715 312
rect 978 441 983 446
rect 811 310 816 315
rect 1044 441 1049 446
rect 979 271 984 276
rect 1068 271 1073 276
rect 729 103 734 108
<< m123contact >>
rect 32 986 37 991
rect 30 955 35 960
rect 32 770 37 775
rect 30 739 35 744
rect 32 554 37 559
rect 30 523 35 528
rect 32 338 37 343
rect 30 307 35 312
rect 32 122 37 127
rect 30 91 35 96
rect 1643 766 1648 771
rect 1641 735 1646 740
rect 1635 466 1640 471
rect 1633 435 1638 440
rect 1635 316 1640 321
rect 1633 285 1638 290
rect 1635 178 1640 183
rect 1633 147 1638 152
<< metal3 >>
rect -20 1010 -13 1011
rect -20 1005 -19 1010
rect -14 1005 -13 1010
rect -20 1004 -13 1005
rect -17 997 -14 1004
rect -9 999 20 1002
rect -9 997 -5 999
rect -17 994 -5 997
rect 17 943 20 999
rect 71 999 78 1000
rect 71 994 72 999
rect 77 994 78 999
rect 71 993 78 994
rect 33 960 36 986
rect 35 957 36 960
rect 17 942 30 943
rect 17 937 24 942
rect 29 937 30 942
rect 17 936 30 937
rect 17 893 20 936
rect 72 897 76 993
rect 805 906 812 907
rect 729 901 806 906
rect 811 901 812 906
rect 81 897 88 898
rect 72 893 82 897
rect 15 892 21 893
rect 81 892 82 893
rect 87 892 88 897
rect 15 887 16 892
rect 21 887 22 892
rect 81 891 88 892
rect 15 886 22 887
rect -20 794 -13 795
rect -20 789 -19 794
rect -14 789 -13 794
rect -20 788 -13 789
rect -17 781 -14 788
rect -9 783 20 786
rect -9 781 -5 783
rect -17 778 -5 781
rect 17 727 20 783
rect 71 783 78 784
rect 71 778 72 783
rect 77 778 78 783
rect 71 777 78 778
rect 33 744 36 770
rect 35 741 36 744
rect 17 726 30 727
rect 17 721 24 726
rect 29 721 30 726
rect 17 720 30 721
rect 17 677 20 720
rect 72 681 76 777
rect 81 681 88 682
rect 72 677 82 681
rect 15 676 21 677
rect 81 676 82 677
rect 87 676 88 681
rect 15 671 16 676
rect 21 671 22 676
rect 81 675 88 676
rect 15 670 22 671
rect -20 578 -13 579
rect -20 573 -19 578
rect -14 573 -13 578
rect -20 572 -13 573
rect -17 565 -14 572
rect -9 567 20 570
rect -9 565 -5 567
rect -17 562 -5 565
rect 17 511 20 567
rect 71 567 78 568
rect 71 562 72 567
rect 77 562 78 567
rect 71 561 78 562
rect 33 528 36 554
rect 35 525 36 528
rect 17 510 30 511
rect 17 505 24 510
rect 29 505 30 510
rect 17 504 30 505
rect 17 461 20 504
rect 72 465 76 561
rect 730 555 734 901
rect 805 900 812 901
rect 1644 740 1647 766
rect 978 739 985 740
rect 978 734 979 739
rect 984 738 985 739
rect 1087 739 1094 740
rect 1087 738 1088 739
rect 984 734 1088 738
rect 1093 734 1094 739
rect 1646 737 1647 740
rect 978 733 985 734
rect 1087 733 1094 734
rect 810 556 817 557
rect 810 555 811 556
rect 730 552 811 555
rect 81 465 88 466
rect 72 461 82 465
rect 15 460 21 461
rect 81 460 82 461
rect 87 460 88 465
rect 15 455 16 460
rect 21 455 22 460
rect 81 459 88 460
rect 15 454 22 455
rect -20 362 -13 363
rect -20 357 -19 362
rect -14 357 -13 362
rect -20 356 -13 357
rect -17 349 -14 356
rect -9 351 20 354
rect -9 349 -5 351
rect -17 346 -5 349
rect 17 295 20 351
rect 71 351 78 352
rect 71 346 72 351
rect 77 346 78 351
rect 71 345 78 346
rect 33 312 36 338
rect 35 309 36 312
rect 17 294 30 295
rect 17 289 24 294
rect 29 289 30 294
rect 17 288 30 289
rect 17 245 20 288
rect 72 249 76 345
rect 730 314 734 552
rect 810 551 811 552
rect 816 551 817 556
rect 810 550 817 551
rect 977 446 984 447
rect 977 441 978 446
rect 983 445 984 446
rect 1043 446 1050 447
rect 1043 445 1044 446
rect 983 441 1044 445
rect 1049 441 1050 446
rect 977 440 984 441
rect 1043 440 1050 441
rect 1636 440 1639 466
rect 1638 437 1639 440
rect 810 315 817 316
rect 810 314 811 315
rect 667 312 674 313
rect 667 307 668 312
rect 673 311 674 312
rect 709 312 716 313
rect 709 311 710 312
rect 673 308 710 311
rect 673 307 674 308
rect 667 306 674 307
rect 709 307 710 308
rect 715 307 716 312
rect 709 306 716 307
rect 730 311 811 314
rect 81 249 88 250
rect 72 245 82 249
rect 15 244 21 245
rect 81 244 82 245
rect 87 244 88 249
rect 15 239 16 244
rect 21 239 22 244
rect 81 243 88 244
rect 15 238 22 239
rect -20 146 -13 147
rect -20 141 -19 146
rect -14 141 -13 146
rect -20 140 -13 141
rect -17 133 -14 140
rect -9 135 20 138
rect -9 133 -5 135
rect -17 130 -5 133
rect 17 79 20 135
rect 71 135 78 136
rect 71 130 72 135
rect 77 130 78 135
rect 71 129 78 130
rect 33 96 36 122
rect 35 93 36 96
rect 17 78 30 79
rect 17 73 24 78
rect 29 73 30 78
rect 17 72 30 73
rect 17 29 20 72
rect 72 33 76 129
rect 730 109 734 311
rect 810 310 811 311
rect 816 310 817 315
rect 810 309 817 310
rect 1636 290 1639 316
rect 1638 287 1639 290
rect 978 276 985 277
rect 978 271 979 276
rect 984 275 985 276
rect 1067 276 1074 277
rect 1067 275 1068 276
rect 984 271 1068 275
rect 1073 271 1074 276
rect 978 270 985 271
rect 1067 270 1074 271
rect 1636 152 1639 178
rect 1638 149 1639 152
rect 728 108 735 109
rect 728 103 729 108
rect 734 103 735 108
rect 728 102 735 103
rect 81 33 88 34
rect 72 29 82 33
rect 15 28 21 29
rect 81 28 82 29
rect 87 28 88 33
rect 15 23 16 28
rect 21 23 22 28
rect 81 27 88 28
rect 15 22 22 23
<< labels >>
rlabel metal1 20 877 20 877 3 gnd
rlabel metal1 20 661 20 661 3 gnd
rlabel metal1 20 445 20 445 3 gnd
rlabel metal1 20 229 20 229 3 gnd
rlabel metal1 20 13 20 13 3 gnd
rlabel metal1 78 878 78 878 7 vdd
rlabel metal1 78 662 78 662 7 vdd
rlabel metal1 78 446 78 446 7 vdd
rlabel metal1 78 230 78 230 7 vdd
rlabel metal1 78 14 78 14 7 vdd
rlabel metal1 2 906 10 910 3 input_1
port 1 s
rlabel metal1 2 690 10 694 3 input_2
port 1 s
rlabel metal1 2 474 10 478 3 input_3
port 1 s
rlabel metal1 2 258 10 262 3 input_4
port 1 s
rlabel metal1 2 42 10 46 3 input_5
port 1 s
rlabel metal1 2 914 10 918 3 input_2
port 2 s
rlabel metal1 2 698 10 702 3 input_3
port 2 s
rlabel metal1 2 482 10 486 3 input_4
port 2 s
rlabel metal1 2 266 10 270 3 input_5
port 2 s
rlabel metal1 2 50 10 54 3 input_6
port 2 s
rlabel metal1 77 918 81 927 7 ground
port 5 n
rlabel metal1 77 702 81 711 7 ground
port 5 n
rlabel metal1 77 486 81 495 7 ground
port 5 n
rlabel metal1 77 270 81 279 7 ground
port 5 n
rlabel metal1 77 54 81 63 7 ground
port 5 n
rlabel metal1 14 919 18 928 5 power_supply
port 3 w
rlabel metal1 14 703 18 712 5 power_supply
port 3 w
rlabel metal1 14 487 18 496 5 power_supply
port 3 w
rlabel metal1 14 271 18 280 5 power_supply
port 3 w
rlabel metal1 14 55 18 64 5 power_supply
port 3 w
rlabel metal1 49 898 53 902 1 output
port 4 e
rlabel metal1 49 682 53 686 1 output
port 4 e
rlabel metal1 49 466 53 470 1 output
port 4 e
rlabel metal1 49 250 53 254 1 output
port 4 e
rlabel metal1 49 34 53 38 1 output
port 4 e
rlabel metal1 74 1013 74 1013 7 vdd
rlabel metal1 74 797 74 797 7 vdd
rlabel metal1 74 581 74 581 7 vdd
rlabel metal1 74 365 74 365 7 vdd
rlabel metal1 74 149 74 149 7 vdd
rlabel metal1 34 994 36 997 1 in1
rlabel metal1 34 778 36 781 1 in2
rlabel metal1 34 562 36 565 1 in3
rlabel metal1 34 346 36 349 1 in4
rlabel metal1 34 130 36 133 1 in5
rlabel m2contact 16 988 16 988 3 in1_inv
rlabel m2contact 16 772 16 772 3 in2_inv
rlabel m2contact 16 556 16 556 3 in3_inv
rlabel m2contact 16 340 16 340 3 in4_inv
rlabel m2contact 16 124 16 124 3 in5_inv
rlabel metal3 36 962 36 962 3 in2
rlabel metal3 36 746 36 746 3 in3
rlabel metal3 36 530 36 530 3 in4
rlabel metal3 36 314 36 314 3 in5
rlabel metal3 36 98 36 98 3 in6
rlabel space 432 72 451 98 1 G0
rlabel space 436 115 455 141 1 G1
rlabel space 436 159 455 185 1 P1
rlabel space 435 209 454 235 1 G2
rlabel space 429 315 448 341 1 P2
rlabel space 435 365 454 391 1 G3
rlabel space 427 557 446 583 1 P3
rlabel space 430 626 449 652 1 G4
rlabel space 416 926 435 952 1 P4
rlabel space 1367 74 1396 100 1 C1
rlabel space 1366 156 1395 182 1 C2
rlabel space 1374 288 1403 314 1 C3
rlabel space 1375 461 1404 487 1 C4
rlabel space 1374 757 1403 783 1 C5
rlabel space 406 -20 435 6 1 ground
rlabel space 427 995 456 1021 5 power
rlabel metal1 1640 454 1640 454 3 out
rlabel metal3 1639 442 1639 442 3 in2
rlabel m2contact 1619 468 1619 468 3 in1_inv
rlabel metal1 1637 474 1639 477 1 in1
rlabel metal1 1618 484 1618 484 3 gnd
rlabel metal1 1677 493 1677 493 7 vdd
rlabel metal1 1640 304 1640 304 3 out
rlabel metal3 1639 292 1639 292 3 in2
rlabel m2contact 1619 318 1619 318 3 in1_inv
rlabel metal1 1637 324 1639 327 1 in1
rlabel metal1 1618 334 1618 334 3 gnd
rlabel metal1 1677 343 1677 343 7 vdd
rlabel metal1 1640 166 1640 166 3 out
rlabel metal3 1639 154 1639 154 3 in2
rlabel m2contact 1619 180 1619 180 3 in1_inv
rlabel metal1 1637 186 1639 189 1 in1
rlabel metal1 1618 196 1618 196 3 gnd
rlabel metal1 1677 205 1677 205 7 vdd
rlabel metal1 1648 754 1648 754 3 out
rlabel metal3 1647 742 1647 742 3 in2
rlabel m2contact 1627 768 1627 768 3 in1_inv
rlabel metal1 1645 774 1647 777 1 in1
rlabel metal1 1626 784 1626 784 3 gnd
rlabel metal1 1685 793 1685 793 7 vdd
<< end >>
