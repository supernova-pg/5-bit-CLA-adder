magic
tech scmos
timestamp 1764778063
<< nwell >>
rect -205 1000 -63 1032
rect 82 998 114 1059
rect -205 917 -63 949
rect 61 937 93 969
rect 958 933 990 989
rect 87 900 119 925
rect 1963 900 2105 932
rect 939 846 971 894
rect -203 785 -61 817
rect 82 782 114 843
rect 929 759 961 799
rect 1253 794 1285 850
rect 1693 778 1725 839
rect 1967 813 2109 845
rect -203 702 -61 734
rect 61 721 93 753
rect 87 684 119 709
rect 894 693 926 725
rect -204 576 -62 608
rect 82 566 114 627
rect 941 581 973 629
rect -204 493 -62 525
rect 61 505 93 537
rect 931 504 963 544
rect 1247 500 1279 548
rect 87 468 119 493
rect 1685 478 1717 539
rect 1959 516 2101 548
rect 894 441 926 473
rect -210 353 -68 385
rect 82 350 114 411
rect 932 341 964 381
rect 1249 326 1281 366
rect 1685 328 1717 389
rect 1959 369 2101 401
rect -210 270 -68 302
rect 61 289 93 321
rect 895 278 927 310
rect 87 252 119 277
rect 893 195 925 227
rect -223 140 -81 172
rect 82 134 114 195
rect 1209 194 1241 226
rect 1685 190 1717 251
rect 1960 222 2102 254
rect 1960 117 2102 149
rect -223 57 -81 89
rect 61 73 93 105
rect 87 36 119 61
<< ntransistor >>
rect 66 1046 76 1048
rect 65 1018 75 1020
rect 65 1009 75 1011
rect -194 974 -192 994
rect -170 974 -168 994
rect -144 980 -142 990
rect -126 974 -124 994
rect -117 974 -115 994
rect -101 974 -99 994
rect -92 974 -90 994
rect -76 980 -74 990
rect 900 976 950 978
rect 900 968 950 970
rect 900 960 950 962
rect 101 956 121 958
rect 900 952 950 954
rect 101 948 121 950
rect 900 944 950 946
rect -194 891 -192 911
rect -170 891 -168 911
rect -144 897 -142 907
rect -126 891 -124 911
rect -117 891 -115 911
rect -101 891 -99 911
rect -92 891 -90 911
rect 71 912 81 914
rect -76 897 -74 907
rect 893 881 933 883
rect 893 873 933 875
rect 1974 874 1976 894
rect 893 865 933 867
rect 1998 874 2000 894
rect 2024 880 2026 890
rect 2042 874 2044 894
rect 2051 874 2053 894
rect 2067 874 2069 894
rect 2076 874 2078 894
rect 2092 880 2094 890
rect 893 857 933 859
rect 1195 837 1245 839
rect 66 830 76 832
rect 1195 829 1245 831
rect 1677 826 1687 828
rect 1195 821 1245 823
rect 1195 813 1245 815
rect 1195 805 1245 807
rect 65 802 75 804
rect 1676 798 1686 800
rect 65 793 75 795
rect -192 759 -190 779
rect -168 759 -166 779
rect -142 765 -140 775
rect -124 759 -122 779
rect -115 759 -113 779
rect -99 759 -97 779
rect -90 759 -88 779
rect 1676 789 1686 791
rect 888 786 918 788
rect 1978 787 1980 807
rect 888 778 918 780
rect 2002 787 2004 807
rect -74 765 -72 775
rect 2028 793 2030 803
rect 2046 787 2048 807
rect 2055 787 2057 807
rect 2071 787 2073 807
rect 2080 787 2082 807
rect 2096 793 2098 803
rect 888 770 918 772
rect 101 740 121 742
rect 101 732 121 734
rect 934 712 954 714
rect -192 676 -190 696
rect -168 676 -166 696
rect -142 682 -140 692
rect -124 676 -122 696
rect -115 676 -113 696
rect -99 676 -97 696
rect -90 676 -88 696
rect 934 704 954 706
rect 71 696 81 698
rect -74 682 -72 692
rect 66 614 76 616
rect 895 616 935 618
rect 895 608 935 610
rect 895 600 935 602
rect 895 592 935 594
rect 65 586 75 588
rect -193 550 -191 570
rect -169 550 -167 570
rect -143 556 -141 566
rect -125 550 -123 570
rect -116 550 -114 570
rect -100 550 -98 570
rect -91 550 -89 570
rect 65 577 75 579
rect -75 556 -73 566
rect 1201 535 1241 537
rect 890 531 920 533
rect 101 524 121 526
rect 1201 527 1241 529
rect 890 523 920 525
rect 101 516 121 518
rect 890 515 920 517
rect 1669 526 1679 528
rect 1201 519 1241 521
rect 1201 511 1241 513
rect -193 467 -191 487
rect -169 467 -167 487
rect -143 473 -141 483
rect -125 467 -123 487
rect -116 467 -114 487
rect -100 467 -98 487
rect -91 467 -89 487
rect 1668 498 1678 500
rect 1668 489 1678 491
rect 1970 490 1972 510
rect -75 473 -73 483
rect 71 480 81 482
rect 1994 490 1996 510
rect 2020 496 2022 506
rect 2038 490 2040 510
rect 2047 490 2049 510
rect 2063 490 2065 510
rect 2072 490 2074 510
rect 2088 496 2090 506
rect 934 460 954 462
rect 934 452 954 454
rect 66 398 76 400
rect 1669 376 1679 378
rect 65 370 75 372
rect 891 368 921 370
rect 65 361 75 363
rect -199 327 -197 347
rect -175 327 -173 347
rect -149 333 -147 343
rect -131 327 -129 347
rect -122 327 -120 347
rect -106 327 -104 347
rect -97 327 -95 347
rect 891 360 921 362
rect 891 352 921 354
rect 1208 353 1238 355
rect 1668 348 1678 350
rect 1208 345 1238 347
rect -81 333 -79 343
rect 1970 343 1972 363
rect 1668 339 1678 341
rect 1208 337 1238 339
rect 1994 343 1996 363
rect 2020 349 2022 359
rect 2038 343 2040 363
rect 2047 343 2049 363
rect 2063 343 2065 363
rect 2072 343 2074 363
rect 2088 349 2090 359
rect 101 308 121 310
rect 101 300 121 302
rect 935 297 955 299
rect 935 289 955 291
rect -199 244 -197 264
rect -175 244 -173 264
rect -149 250 -147 260
rect -131 244 -129 264
rect -122 244 -120 264
rect -106 244 -104 264
rect -97 244 -95 264
rect 71 264 81 266
rect -81 250 -79 260
rect 1669 238 1679 240
rect 933 214 953 216
rect 1249 213 1269 215
rect 933 206 953 208
rect 1668 210 1678 212
rect 1249 205 1269 207
rect 1668 201 1678 203
rect 1971 196 1973 216
rect 1995 196 1997 216
rect 66 182 76 184
rect 2021 202 2023 212
rect 2039 196 2041 216
rect 2048 196 2050 216
rect 2064 196 2066 216
rect 2073 196 2075 216
rect 2089 202 2091 212
rect 65 154 75 156
rect -212 114 -210 134
rect -188 114 -186 134
rect -162 120 -160 130
rect -144 114 -142 134
rect -135 114 -133 134
rect -119 114 -117 134
rect -110 114 -108 134
rect 65 145 75 147
rect -94 120 -92 130
rect 101 92 121 94
rect 1971 91 1973 111
rect 101 84 121 86
rect 1995 91 1997 111
rect 2021 97 2023 107
rect 2039 91 2041 111
rect 2048 91 2050 111
rect 2064 91 2066 111
rect 2073 91 2075 111
rect 2089 97 2091 107
rect -212 31 -210 51
rect -188 31 -186 51
rect -162 37 -160 47
rect -144 31 -142 51
rect -135 31 -133 51
rect -119 31 -117 51
rect -110 31 -108 51
rect 71 48 81 50
rect -94 37 -92 47
<< ptransistor >>
rect 88 1046 108 1048
rect -194 1006 -192 1026
rect -186 1006 -184 1026
rect -170 1006 -168 1026
rect -162 1006 -160 1026
rect -144 1006 -142 1026
rect -126 1006 -124 1026
rect -101 1006 -99 1026
rect -76 1006 -74 1026
rect 88 1018 108 1020
rect 88 1009 108 1011
rect 964 976 984 978
rect 964 968 984 970
rect 964 960 984 962
rect 67 956 87 958
rect 964 952 984 954
rect 67 948 87 950
rect 964 944 984 946
rect -194 923 -192 943
rect -186 923 -184 943
rect -170 923 -168 943
rect -162 923 -160 943
rect -144 923 -142 943
rect -126 923 -124 943
rect -101 923 -99 943
rect -76 923 -74 943
rect 93 912 113 914
rect 1974 906 1976 926
rect 1982 906 1984 926
rect 1998 906 2000 926
rect 2006 906 2008 926
rect 2024 906 2026 926
rect 2042 906 2044 926
rect 2067 906 2069 926
rect 2092 906 2094 926
rect 945 881 965 883
rect 945 873 965 875
rect 945 865 965 867
rect 945 857 965 859
rect 1259 837 1279 839
rect 88 830 108 832
rect 1259 829 1279 831
rect 1699 826 1719 828
rect 1259 821 1279 823
rect 1978 819 1980 839
rect 1986 819 1988 839
rect 2002 819 2004 839
rect 2010 819 2012 839
rect 2028 819 2030 839
rect 2046 819 2048 839
rect 2071 819 2073 839
rect 2096 819 2098 839
rect 1259 813 1279 815
rect -192 791 -190 811
rect -184 791 -182 811
rect -168 791 -166 811
rect -160 791 -158 811
rect -142 791 -140 811
rect -124 791 -122 811
rect -99 791 -97 811
rect -74 791 -72 811
rect 1259 805 1279 807
rect 88 802 108 804
rect 1699 798 1719 800
rect 88 793 108 795
rect 1699 789 1719 791
rect 935 786 955 788
rect 935 778 955 780
rect 935 770 955 772
rect 67 740 87 742
rect 67 732 87 734
rect -192 708 -190 728
rect -184 708 -182 728
rect -168 708 -166 728
rect -160 708 -158 728
rect -142 708 -140 728
rect -124 708 -122 728
rect -99 708 -97 728
rect -74 708 -72 728
rect 900 712 920 714
rect 900 704 920 706
rect 93 696 113 698
rect 88 614 108 616
rect 947 616 967 618
rect 947 608 967 610
rect -193 582 -191 602
rect -185 582 -183 602
rect -169 582 -167 602
rect -161 582 -159 602
rect -143 582 -141 602
rect -125 582 -123 602
rect -100 582 -98 602
rect -75 582 -73 602
rect 947 600 967 602
rect 947 592 967 594
rect 88 586 108 588
rect 88 577 108 579
rect 1253 535 1273 537
rect 937 531 957 533
rect 67 524 87 526
rect -193 499 -191 519
rect -185 499 -183 519
rect -169 499 -167 519
rect -161 499 -159 519
rect -143 499 -141 519
rect -125 499 -123 519
rect -100 499 -98 519
rect -75 499 -73 519
rect 1253 527 1273 529
rect 937 523 957 525
rect 67 516 87 518
rect 937 515 957 517
rect 1691 526 1711 528
rect 1970 522 1972 542
rect 1978 522 1980 542
rect 1994 522 1996 542
rect 2002 522 2004 542
rect 2020 522 2022 542
rect 2038 522 2040 542
rect 2063 522 2065 542
rect 2088 522 2090 542
rect 1253 519 1273 521
rect 1253 511 1273 513
rect 1691 498 1711 500
rect 1691 489 1711 491
rect 93 480 113 482
rect 900 460 920 462
rect 900 452 920 454
rect 88 398 108 400
rect -199 359 -197 379
rect -191 359 -189 379
rect -175 359 -173 379
rect -167 359 -165 379
rect -149 359 -147 379
rect -131 359 -129 379
rect -106 359 -104 379
rect -81 359 -79 379
rect 1691 376 1711 378
rect 88 370 108 372
rect 1970 375 1972 395
rect 1978 375 1980 395
rect 1994 375 1996 395
rect 2002 375 2004 395
rect 2020 375 2022 395
rect 2038 375 2040 395
rect 2063 375 2065 395
rect 2088 375 2090 395
rect 938 368 958 370
rect 88 361 108 363
rect 938 360 958 362
rect 938 352 958 354
rect 1255 353 1275 355
rect 1691 348 1711 350
rect 1255 345 1275 347
rect 1691 339 1711 341
rect 1255 337 1275 339
rect 67 308 87 310
rect 67 300 87 302
rect -199 276 -197 296
rect -191 276 -189 296
rect -175 276 -173 296
rect -167 276 -165 296
rect -149 276 -147 296
rect -131 276 -129 296
rect -106 276 -104 296
rect -81 276 -79 296
rect 901 297 921 299
rect 901 289 921 291
rect 93 264 113 266
rect 1691 238 1711 240
rect 1971 228 1973 248
rect 1979 228 1981 248
rect 1995 228 1997 248
rect 2003 228 2005 248
rect 2021 228 2023 248
rect 2039 228 2041 248
rect 2064 228 2066 248
rect 2089 228 2091 248
rect 899 214 919 216
rect 1215 213 1235 215
rect 899 206 919 208
rect 1691 210 1711 212
rect 1215 205 1235 207
rect 1691 201 1711 203
rect 88 182 108 184
rect -212 146 -210 166
rect -204 146 -202 166
rect -188 146 -186 166
rect -180 146 -178 166
rect -162 146 -160 166
rect -144 146 -142 166
rect -119 146 -117 166
rect -94 146 -92 166
rect 88 154 108 156
rect 88 145 108 147
rect 1971 123 1973 143
rect 1979 123 1981 143
rect 1995 123 1997 143
rect 2003 123 2005 143
rect 2021 123 2023 143
rect 2039 123 2041 143
rect 2064 123 2066 143
rect 2089 123 2091 143
rect 67 92 87 94
rect 67 84 87 86
rect -212 63 -210 83
rect -204 63 -202 83
rect -188 63 -186 83
rect -180 63 -178 83
rect -162 63 -160 83
rect -144 63 -142 83
rect -119 63 -117 83
rect -94 63 -92 83
rect 93 48 113 50
<< ndiffusion >>
rect 70 1049 76 1053
rect 66 1048 76 1049
rect 66 1045 76 1046
rect 70 1041 76 1045
rect 69 1021 75 1025
rect 65 1020 75 1021
rect 65 1017 75 1018
rect 65 1013 71 1017
rect 65 1011 75 1013
rect 65 1008 75 1009
rect -199 978 -194 994
rect -195 974 -194 978
rect -192 990 -191 994
rect -192 974 -187 990
rect -175 978 -170 994
rect -171 974 -170 978
rect -168 990 -167 994
rect -168 974 -163 990
rect -149 984 -144 990
rect -145 980 -144 984
rect -142 986 -141 990
rect -142 980 -137 986
rect -131 978 -126 994
rect -127 974 -126 978
rect -124 974 -117 994
rect -115 990 -114 994
rect -115 974 -110 990
rect -106 978 -101 994
rect -102 974 -101 978
rect -99 974 -92 994
rect -90 990 -89 994
rect 65 1004 71 1008
rect -90 974 -85 990
rect -81 984 -76 990
rect -77 980 -76 984
rect -74 986 -73 990
rect -74 980 -69 986
rect 900 978 950 979
rect 900 975 950 976
rect 900 970 950 971
rect 900 967 950 968
rect 900 962 950 963
rect 900 959 950 960
rect 101 958 121 959
rect 101 955 121 956
rect 900 954 950 955
rect 900 951 950 952
rect 101 950 121 951
rect 101 947 121 948
rect 900 946 950 947
rect 900 943 950 944
rect -199 895 -194 911
rect -195 891 -194 895
rect -192 907 -191 911
rect -192 891 -187 907
rect -175 895 -170 911
rect -171 891 -170 895
rect -168 907 -167 911
rect -168 891 -163 907
rect -149 901 -144 907
rect -145 897 -144 901
rect -142 903 -141 907
rect -142 897 -137 903
rect -131 895 -126 911
rect -127 891 -126 895
rect -124 891 -117 911
rect -115 907 -114 911
rect -115 891 -110 907
rect -106 895 -101 911
rect -102 891 -101 895
rect -99 891 -92 911
rect -90 907 -89 911
rect 75 915 81 919
rect 71 914 81 915
rect 71 911 81 912
rect 71 907 77 911
rect -90 891 -85 907
rect -81 901 -76 907
rect -77 897 -76 901
rect -74 903 -73 907
rect -74 897 -69 903
rect 893 883 933 884
rect 893 880 933 881
rect 893 875 933 876
rect 1969 878 1974 894
rect 1973 874 1974 878
rect 1976 890 1977 894
rect 1976 874 1981 890
rect 893 872 933 873
rect 893 867 933 868
rect 1993 878 1998 894
rect 1997 874 1998 878
rect 2000 890 2001 894
rect 2000 874 2005 890
rect 893 864 933 865
rect 893 859 933 860
rect 2019 884 2024 890
rect 2023 880 2024 884
rect 2026 886 2027 890
rect 2026 880 2031 886
rect 2037 878 2042 894
rect 2041 874 2042 878
rect 2044 874 2051 894
rect 2053 890 2054 894
rect 2053 874 2058 890
rect 2062 878 2067 894
rect 2066 874 2067 878
rect 2069 874 2076 894
rect 2078 890 2079 894
rect 2078 874 2083 890
rect 2087 884 2092 890
rect 2091 880 2092 884
rect 2094 886 2095 890
rect 2094 880 2099 886
rect 893 856 933 857
rect 70 833 76 837
rect 66 832 76 833
rect 1195 839 1245 840
rect 1195 836 1245 837
rect 66 829 76 830
rect 70 825 76 829
rect 1195 831 1245 832
rect 1681 829 1687 833
rect 1195 828 1245 829
rect 1195 823 1245 824
rect 1677 828 1687 829
rect 1677 825 1687 826
rect 1681 821 1687 825
rect 1195 820 1245 821
rect 1195 815 1245 816
rect 1195 812 1245 813
rect 69 805 75 809
rect 65 804 75 805
rect 1195 807 1245 808
rect 1195 804 1245 805
rect 65 801 75 802
rect 65 797 71 801
rect 65 795 75 797
rect 1680 801 1686 805
rect 1676 800 1686 801
rect 1676 797 1686 798
rect 65 792 75 793
rect -197 763 -192 779
rect -193 759 -192 763
rect -190 775 -189 779
rect -190 759 -185 775
rect -173 763 -168 779
rect -169 759 -168 763
rect -166 775 -165 779
rect -166 759 -161 775
rect -147 769 -142 775
rect -143 765 -142 769
rect -140 771 -139 775
rect -140 765 -135 771
rect -129 763 -124 779
rect -125 759 -124 763
rect -122 759 -115 779
rect -113 775 -112 779
rect -113 759 -108 775
rect -104 763 -99 779
rect -100 759 -99 763
rect -97 759 -90 779
rect -88 775 -87 779
rect 65 788 71 792
rect 888 788 918 789
rect 1676 793 1682 797
rect 1676 791 1686 793
rect 1973 791 1978 807
rect 1676 788 1686 789
rect 888 785 918 786
rect 888 780 918 781
rect 1676 784 1682 788
rect 1977 787 1978 791
rect 1980 803 1981 807
rect 1980 787 1985 803
rect 1997 791 2002 807
rect 2001 787 2002 791
rect 2004 803 2005 807
rect 2004 787 2009 803
rect 888 777 918 778
rect -88 759 -83 775
rect -79 769 -74 775
rect -75 765 -74 769
rect -72 771 -71 775
rect -72 765 -67 771
rect 888 772 918 773
rect 2023 797 2028 803
rect 2027 793 2028 797
rect 2030 799 2031 803
rect 2030 793 2035 799
rect 2041 791 2046 807
rect 2045 787 2046 791
rect 2048 787 2055 807
rect 2057 803 2058 807
rect 2057 787 2062 803
rect 2066 791 2071 807
rect 2070 787 2071 791
rect 2073 787 2080 807
rect 2082 803 2083 807
rect 2082 787 2087 803
rect 2091 797 2096 803
rect 2095 793 2096 797
rect 2098 799 2099 803
rect 2098 793 2103 799
rect 888 769 918 770
rect 101 742 121 743
rect 101 739 121 740
rect 101 734 121 735
rect 101 731 121 732
rect 934 714 954 715
rect -197 680 -192 696
rect -193 676 -192 680
rect -190 692 -189 696
rect -190 676 -185 692
rect -173 680 -168 696
rect -169 676 -168 680
rect -166 692 -165 696
rect -166 676 -161 692
rect -147 686 -142 692
rect -143 682 -142 686
rect -140 688 -139 692
rect -140 682 -135 688
rect -129 680 -124 696
rect -125 676 -124 680
rect -122 676 -115 696
rect -113 692 -112 696
rect -113 676 -108 692
rect -104 680 -99 696
rect -100 676 -99 680
rect -97 676 -90 696
rect -88 692 -87 696
rect 934 711 954 712
rect 934 706 954 707
rect 75 699 81 703
rect 71 698 81 699
rect 934 703 954 704
rect 71 695 81 696
rect -88 676 -83 692
rect -79 686 -74 692
rect -75 682 -74 686
rect -72 688 -71 692
rect 71 691 77 695
rect -72 682 -67 688
rect 70 617 76 621
rect 66 616 76 617
rect 895 618 935 619
rect 895 615 935 616
rect 66 613 76 614
rect 70 609 76 613
rect 895 610 935 611
rect 895 607 935 608
rect 895 602 935 603
rect 895 599 935 600
rect 69 589 75 593
rect 65 588 75 589
rect 895 594 935 595
rect 895 591 935 592
rect 65 585 75 586
rect -198 554 -193 570
rect -194 550 -193 554
rect -191 566 -190 570
rect -191 550 -186 566
rect -174 554 -169 570
rect -170 550 -169 554
rect -167 566 -166 570
rect -167 550 -162 566
rect -148 560 -143 566
rect -144 556 -143 560
rect -141 562 -140 566
rect -141 556 -136 562
rect -130 554 -125 570
rect -126 550 -125 554
rect -123 550 -116 570
rect -114 566 -113 570
rect -114 550 -109 566
rect -105 554 -100 570
rect -101 550 -100 554
rect -98 550 -91 570
rect -89 566 -88 570
rect 65 581 71 585
rect 65 579 75 581
rect 65 576 75 577
rect 65 572 71 576
rect -89 550 -84 566
rect -80 560 -75 566
rect -76 556 -75 560
rect -73 562 -72 566
rect -73 556 -68 562
rect 890 533 920 534
rect 1201 537 1241 538
rect 1201 534 1241 535
rect 890 530 920 531
rect 101 526 121 527
rect 101 523 121 524
rect 890 525 920 526
rect 1201 529 1241 530
rect 1673 529 1679 533
rect 1669 528 1679 529
rect 1201 526 1241 527
rect 890 522 920 523
rect 101 518 121 519
rect 101 515 121 516
rect 890 517 920 518
rect 890 514 920 515
rect 1201 521 1241 522
rect 1669 525 1679 526
rect 1673 521 1679 525
rect 1201 518 1241 519
rect 1201 513 1241 514
rect 1201 510 1241 511
rect 1672 501 1678 505
rect 1668 500 1678 501
rect -198 471 -193 487
rect -194 467 -193 471
rect -191 483 -190 487
rect -191 467 -186 483
rect -174 471 -169 487
rect -170 467 -169 471
rect -167 483 -166 487
rect -167 467 -162 483
rect -148 477 -143 483
rect -144 473 -143 477
rect -141 479 -140 483
rect -141 473 -136 479
rect -130 471 -125 487
rect -126 467 -125 471
rect -123 467 -116 487
rect -114 483 -113 487
rect -114 467 -109 483
rect -105 471 -100 487
rect -101 467 -100 471
rect -98 467 -91 487
rect -89 483 -88 487
rect 1668 497 1678 498
rect 1668 493 1674 497
rect 1668 491 1678 493
rect 1965 494 1970 510
rect 1969 490 1970 494
rect 1972 506 1973 510
rect 1972 490 1977 506
rect 1668 488 1678 489
rect 75 483 81 487
rect -89 467 -84 483
rect -80 477 -75 483
rect -76 473 -75 477
rect -73 479 -72 483
rect 71 482 81 483
rect 1668 484 1674 488
rect 1989 494 1994 510
rect 1993 490 1994 494
rect 1996 506 1997 510
rect 1996 490 2001 506
rect -73 473 -68 479
rect 71 479 81 480
rect 71 475 77 479
rect 2015 500 2020 506
rect 2019 496 2020 500
rect 2022 502 2023 506
rect 2022 496 2027 502
rect 2033 494 2038 510
rect 2037 490 2038 494
rect 2040 490 2047 510
rect 2049 506 2050 510
rect 2049 490 2054 506
rect 2058 494 2063 510
rect 2062 490 2063 494
rect 2065 490 2072 510
rect 2074 506 2075 510
rect 2074 490 2079 506
rect 2083 500 2088 506
rect 2087 496 2088 500
rect 2090 502 2091 506
rect 2090 496 2095 502
rect 934 462 954 463
rect 934 459 954 460
rect 934 454 954 455
rect 934 451 954 452
rect 70 401 76 405
rect 66 400 76 401
rect 66 397 76 398
rect 70 393 76 397
rect 1673 379 1679 383
rect 1669 378 1679 379
rect 69 373 75 377
rect 65 372 75 373
rect 1669 375 1679 376
rect 65 369 75 370
rect 65 365 71 369
rect 65 363 75 365
rect 891 370 921 371
rect 1673 371 1679 375
rect 891 367 921 368
rect 65 360 75 361
rect -204 331 -199 347
rect -200 327 -199 331
rect -197 343 -196 347
rect -197 327 -192 343
rect -180 331 -175 347
rect -176 327 -175 331
rect -173 343 -172 347
rect -173 327 -168 343
rect -154 337 -149 343
rect -150 333 -149 337
rect -147 339 -146 343
rect -147 333 -142 339
rect -136 331 -131 347
rect -132 327 -131 331
rect -129 327 -122 347
rect -120 343 -119 347
rect -120 327 -115 343
rect -111 331 -106 347
rect -107 327 -106 331
rect -104 327 -97 347
rect -95 343 -94 347
rect 65 356 71 360
rect 891 362 921 363
rect 891 359 921 360
rect 891 354 921 355
rect 1208 355 1238 356
rect 1208 352 1238 353
rect 891 351 921 352
rect 1208 347 1238 348
rect 1672 351 1678 355
rect 1668 350 1678 351
rect 1668 347 1678 348
rect 1208 344 1238 345
rect -95 327 -90 343
rect -86 337 -81 343
rect -82 333 -81 337
rect -79 339 -78 343
rect -79 333 -74 339
rect 1208 339 1238 340
rect 1668 343 1674 347
rect 1668 341 1678 343
rect 1965 347 1970 363
rect 1969 343 1970 347
rect 1972 359 1973 363
rect 1972 343 1977 359
rect 1668 338 1678 339
rect 1208 336 1238 337
rect 1668 334 1674 338
rect 1989 347 1994 363
rect 1993 343 1994 347
rect 1996 359 1997 363
rect 1996 343 2001 359
rect 2015 353 2020 359
rect 2019 349 2020 353
rect 2022 355 2023 359
rect 2022 349 2027 355
rect 2033 347 2038 363
rect 2037 343 2038 347
rect 2040 343 2047 363
rect 2049 359 2050 363
rect 2049 343 2054 359
rect 2058 347 2063 363
rect 2062 343 2063 347
rect 2065 343 2072 363
rect 2074 359 2075 363
rect 2074 343 2079 359
rect 2083 353 2088 359
rect 2087 349 2088 353
rect 2090 355 2091 359
rect 2090 349 2095 355
rect 101 310 121 311
rect 101 307 121 308
rect 101 302 121 303
rect 101 299 121 300
rect 935 299 955 300
rect 935 296 955 297
rect 935 291 955 292
rect 935 288 955 289
rect -204 248 -199 264
rect -200 244 -199 248
rect -197 260 -196 264
rect -197 244 -192 260
rect -180 248 -175 264
rect -176 244 -175 248
rect -173 260 -172 264
rect -173 244 -168 260
rect -154 254 -149 260
rect -150 250 -149 254
rect -147 256 -146 260
rect -147 250 -142 256
rect -136 248 -131 264
rect -132 244 -131 248
rect -129 244 -122 264
rect -120 260 -119 264
rect -120 244 -115 260
rect -111 248 -106 264
rect -107 244 -106 248
rect -104 244 -97 264
rect -95 260 -94 264
rect 75 267 81 271
rect 71 266 81 267
rect 71 263 81 264
rect -95 244 -90 260
rect -86 254 -81 260
rect -82 250 -81 254
rect -79 256 -78 260
rect 71 259 77 263
rect -79 250 -74 256
rect 1673 241 1679 245
rect 1669 240 1679 241
rect 1669 237 1679 238
rect 1673 233 1679 237
rect 933 216 953 217
rect 933 213 953 214
rect 1249 215 1269 216
rect 1672 213 1678 217
rect 933 208 953 209
rect 933 205 953 206
rect 1249 212 1269 213
rect 1668 212 1678 213
rect 1249 207 1269 208
rect 1668 209 1678 210
rect 1249 204 1269 205
rect 1668 205 1674 209
rect 1668 203 1678 205
rect 1668 200 1678 201
rect 1668 196 1674 200
rect 1966 200 1971 216
rect 1970 196 1971 200
rect 1973 212 1974 216
rect 1973 196 1978 212
rect 70 185 76 189
rect 66 184 76 185
rect 1990 200 1995 216
rect 1994 196 1995 200
rect 1997 212 1998 216
rect 1997 196 2002 212
rect 2016 206 2021 212
rect 2020 202 2021 206
rect 2023 208 2024 212
rect 2023 202 2028 208
rect 2034 200 2039 216
rect 2038 196 2039 200
rect 2041 196 2048 216
rect 2050 212 2051 216
rect 2050 196 2055 212
rect 2059 200 2064 216
rect 2063 196 2064 200
rect 2066 196 2073 216
rect 2075 212 2076 216
rect 2075 196 2080 212
rect 2084 206 2089 212
rect 2088 202 2089 206
rect 2091 208 2092 212
rect 2091 202 2096 208
rect 66 181 76 182
rect 70 177 76 181
rect 69 157 75 161
rect 65 156 75 157
rect 65 153 75 154
rect 65 149 71 153
rect 65 147 75 149
rect -217 118 -212 134
rect -213 114 -212 118
rect -210 130 -209 134
rect -210 114 -205 130
rect -193 118 -188 134
rect -189 114 -188 118
rect -186 130 -185 134
rect -186 114 -181 130
rect -167 124 -162 130
rect -163 120 -162 124
rect -160 126 -159 130
rect -160 120 -155 126
rect -149 118 -144 134
rect -145 114 -144 118
rect -142 114 -135 134
rect -133 130 -132 134
rect -133 114 -128 130
rect -124 118 -119 134
rect -120 114 -119 118
rect -117 114 -110 134
rect -108 130 -107 134
rect 65 144 75 145
rect 65 140 71 144
rect -108 114 -103 130
rect -99 124 -94 130
rect -95 120 -94 124
rect -92 126 -91 130
rect -92 120 -87 126
rect 101 94 121 95
rect 1966 95 1971 111
rect 101 91 121 92
rect 1970 91 1971 95
rect 1973 107 1974 111
rect 1973 91 1978 107
rect 101 86 121 87
rect 101 83 121 84
rect 1990 95 1995 111
rect 1994 91 1995 95
rect 1997 107 1998 111
rect 1997 91 2002 107
rect 2016 101 2021 107
rect 2020 97 2021 101
rect 2023 103 2024 107
rect 2023 97 2028 103
rect 2034 95 2039 111
rect 2038 91 2039 95
rect 2041 91 2048 111
rect 2050 107 2051 111
rect 2050 91 2055 107
rect 2059 95 2064 111
rect 2063 91 2064 95
rect 2066 91 2073 111
rect 2075 107 2076 111
rect 2075 91 2080 107
rect 2084 101 2089 107
rect 2088 97 2089 101
rect 2091 103 2092 107
rect 2091 97 2096 103
rect -217 35 -212 51
rect -213 31 -212 35
rect -210 47 -209 51
rect -210 31 -205 47
rect -193 35 -188 51
rect -189 31 -188 35
rect -186 47 -185 51
rect -186 31 -181 47
rect -167 41 -162 47
rect -163 37 -162 41
rect -160 43 -159 47
rect -160 37 -155 43
rect -149 35 -144 51
rect -145 31 -144 35
rect -142 31 -135 51
rect -133 47 -132 51
rect -133 31 -128 47
rect -124 35 -119 51
rect -120 31 -119 35
rect -117 31 -110 51
rect -108 47 -107 51
rect 75 51 81 55
rect 71 50 81 51
rect 71 47 81 48
rect -108 31 -103 47
rect -99 41 -94 47
rect -95 37 -94 41
rect -92 43 -91 47
rect 71 43 77 47
rect -92 37 -87 43
<< pdiffusion >>
rect 92 1049 108 1053
rect 88 1048 108 1049
rect 88 1045 108 1046
rect 88 1041 104 1045
rect -195 1022 -194 1026
rect -199 1006 -194 1022
rect -192 1006 -186 1026
rect -184 1010 -179 1026
rect -184 1006 -183 1010
rect -171 1022 -170 1026
rect -175 1006 -170 1022
rect -168 1006 -162 1026
rect -160 1010 -155 1026
rect -160 1006 -159 1010
rect -145 1022 -144 1026
rect -149 1006 -144 1022
rect -142 1010 -137 1026
rect -142 1006 -141 1010
rect -127 1022 -126 1026
rect -131 1006 -126 1022
rect -124 1010 -119 1026
rect -124 1006 -123 1010
rect -102 1022 -101 1026
rect -106 1006 -101 1022
rect -99 1010 -94 1026
rect -99 1006 -98 1010
rect -77 1022 -76 1026
rect -81 1006 -76 1022
rect -74 1010 -69 1026
rect 88 1021 104 1025
rect 88 1020 108 1021
rect -74 1006 -73 1010
rect 88 1017 108 1018
rect 88 1013 90 1017
rect 94 1013 108 1017
rect 88 1011 108 1013
rect 88 1008 108 1009
rect 92 1004 108 1008
rect 964 978 984 979
rect 964 975 984 976
rect 964 970 984 971
rect 67 958 87 959
rect 964 967 984 968
rect 964 962 984 963
rect 67 955 87 956
rect 67 950 87 951
rect 964 959 984 960
rect 964 954 984 955
rect 67 947 87 948
rect 964 951 984 952
rect 964 946 984 947
rect -195 939 -194 943
rect -199 923 -194 939
rect -192 923 -186 943
rect -184 927 -179 943
rect -184 923 -183 927
rect -171 939 -170 943
rect -175 923 -170 939
rect -168 923 -162 943
rect -160 927 -155 943
rect -160 923 -159 927
rect -145 939 -144 943
rect -149 923 -144 939
rect -142 927 -137 943
rect -142 923 -141 927
rect -127 939 -126 943
rect -131 923 -126 939
rect -124 927 -119 943
rect -124 923 -123 927
rect -102 939 -101 943
rect -106 923 -101 939
rect -99 927 -94 943
rect -99 923 -98 927
rect -77 939 -76 943
rect -81 923 -76 939
rect -74 927 -69 943
rect 964 943 984 944
rect -74 923 -73 927
rect 1973 922 1974 926
rect 93 915 109 919
rect 93 914 113 915
rect 93 911 113 912
rect 97 907 113 911
rect 1969 906 1974 922
rect 1976 906 1982 926
rect 1984 910 1989 926
rect 1984 906 1985 910
rect 1997 922 1998 926
rect 1993 906 1998 922
rect 2000 906 2006 926
rect 2008 910 2013 926
rect 2008 906 2009 910
rect 2023 922 2024 926
rect 2019 906 2024 922
rect 2026 910 2031 926
rect 2026 906 2027 910
rect 2041 922 2042 926
rect 2037 906 2042 922
rect 2044 910 2049 926
rect 2044 906 2045 910
rect 2066 922 2067 926
rect 2062 906 2067 922
rect 2069 910 2074 926
rect 2069 906 2070 910
rect 2091 922 2092 926
rect 2087 906 2092 922
rect 2094 910 2099 926
rect 2094 906 2095 910
rect 945 883 965 884
rect 945 880 965 881
rect 945 875 965 876
rect 945 872 965 873
rect 945 867 965 868
rect 945 864 965 865
rect 945 859 965 860
rect 945 856 965 857
rect 92 833 108 837
rect 1259 839 1279 840
rect 88 832 108 833
rect 88 829 108 830
rect 88 825 104 829
rect 1259 836 1279 837
rect 1977 835 1978 839
rect 1259 831 1279 832
rect 1259 828 1279 829
rect 1703 829 1719 833
rect 1699 828 1719 829
rect 1259 823 1279 824
rect 1699 825 1719 826
rect 1699 821 1715 825
rect 1259 820 1279 821
rect 1973 819 1978 835
rect 1980 819 1986 839
rect 1988 823 1993 839
rect 1988 819 1989 823
rect 2001 835 2002 839
rect 1997 819 2002 835
rect 2004 819 2010 839
rect 2012 823 2017 839
rect 2012 819 2013 823
rect 2027 835 2028 839
rect 2023 819 2028 835
rect 2030 823 2035 839
rect 2030 819 2031 823
rect 2045 835 2046 839
rect 2041 819 2046 835
rect 2048 823 2053 839
rect 2048 819 2049 823
rect 2070 835 2071 839
rect 2066 819 2071 835
rect 2073 823 2078 839
rect 2073 819 2074 823
rect 2095 835 2096 839
rect 2091 819 2096 835
rect 2098 823 2103 839
rect 2098 819 2099 823
rect 1259 815 1279 816
rect -193 807 -192 811
rect -197 791 -192 807
rect -190 791 -184 811
rect -182 795 -177 811
rect -182 791 -181 795
rect -169 807 -168 811
rect -173 791 -168 807
rect -166 791 -160 811
rect -158 795 -153 811
rect -158 791 -157 795
rect -143 807 -142 811
rect -147 791 -142 807
rect -140 795 -135 811
rect -140 791 -139 795
rect -125 807 -124 811
rect -129 791 -124 807
rect -122 795 -117 811
rect -122 791 -121 795
rect -100 807 -99 811
rect -104 791 -99 807
rect -97 795 -92 811
rect -97 791 -96 795
rect -75 807 -74 811
rect -79 791 -74 807
rect -72 795 -67 811
rect 88 805 104 809
rect 88 804 108 805
rect 1259 812 1279 813
rect 1259 807 1279 808
rect -72 791 -71 795
rect 88 801 108 802
rect 88 797 90 801
rect 94 797 108 801
rect 1259 804 1279 805
rect 1699 801 1715 805
rect 1699 800 1719 801
rect 88 795 108 797
rect 88 792 108 793
rect 92 788 108 792
rect 1699 797 1719 798
rect 1699 793 1701 797
rect 1705 793 1719 797
rect 1699 791 1719 793
rect 935 788 955 789
rect 935 785 955 786
rect 1699 788 1719 789
rect 1703 784 1719 788
rect 935 780 955 781
rect 935 777 955 778
rect 935 772 955 773
rect 935 769 955 770
rect 67 742 87 743
rect 67 739 87 740
rect 67 734 87 735
rect 67 731 87 732
rect -193 724 -192 728
rect -197 708 -192 724
rect -190 708 -184 728
rect -182 712 -177 728
rect -182 708 -181 712
rect -169 724 -168 728
rect -173 708 -168 724
rect -166 708 -160 728
rect -158 712 -153 728
rect -158 708 -157 712
rect -143 724 -142 728
rect -147 708 -142 724
rect -140 712 -135 728
rect -140 708 -139 712
rect -125 724 -124 728
rect -129 708 -124 724
rect -122 712 -117 728
rect -122 708 -121 712
rect -100 724 -99 728
rect -104 708 -99 724
rect -97 712 -92 728
rect -97 708 -96 712
rect -75 724 -74 728
rect -79 708 -74 724
rect -72 712 -67 728
rect -72 708 -71 712
rect 900 714 920 715
rect 900 711 920 712
rect 900 706 920 707
rect 900 703 920 704
rect 93 699 109 703
rect 93 698 113 699
rect 93 695 113 696
rect 97 691 113 695
rect 92 617 108 621
rect 88 616 108 617
rect 947 618 967 619
rect 88 613 108 614
rect 88 609 104 613
rect 947 615 967 616
rect 947 610 967 611
rect -194 598 -193 602
rect -198 582 -193 598
rect -191 582 -185 602
rect -183 586 -178 602
rect -183 582 -182 586
rect -170 598 -169 602
rect -174 582 -169 598
rect -167 582 -161 602
rect -159 586 -154 602
rect -159 582 -158 586
rect -144 598 -143 602
rect -148 582 -143 598
rect -141 586 -136 602
rect -141 582 -140 586
rect -126 598 -125 602
rect -130 582 -125 598
rect -123 586 -118 602
rect -123 582 -122 586
rect -101 598 -100 602
rect -105 582 -100 598
rect -98 586 -93 602
rect -98 582 -97 586
rect -76 598 -75 602
rect -80 582 -75 598
rect -73 586 -68 602
rect 947 607 967 608
rect 947 602 967 603
rect 88 589 104 593
rect 947 599 967 600
rect 947 594 967 595
rect 88 588 108 589
rect 947 591 967 592
rect -73 582 -72 586
rect 88 585 108 586
rect 88 581 90 585
rect 94 581 108 585
rect 88 579 108 581
rect 88 576 108 577
rect 92 572 108 576
rect 67 526 87 527
rect 1253 537 1273 538
rect 1969 538 1970 542
rect 937 533 957 534
rect 67 523 87 524
rect -194 515 -193 519
rect -198 499 -193 515
rect -191 499 -185 519
rect -183 503 -178 519
rect -183 499 -182 503
rect -170 515 -169 519
rect -174 499 -169 515
rect -167 499 -161 519
rect -159 503 -154 519
rect -159 499 -158 503
rect -144 515 -143 519
rect -148 499 -143 515
rect -141 503 -136 519
rect -141 499 -140 503
rect -126 515 -125 519
rect -130 499 -125 515
rect -123 503 -118 519
rect -123 499 -122 503
rect -101 515 -100 519
rect -105 499 -100 515
rect -98 503 -93 519
rect -98 499 -97 503
rect -76 515 -75 519
rect -80 499 -75 515
rect -73 503 -68 519
rect 67 518 87 519
rect 937 530 957 531
rect 1253 534 1273 535
rect 1253 529 1273 530
rect 1695 529 1711 533
rect 1691 528 1711 529
rect 937 525 957 526
rect 67 515 87 516
rect 937 522 957 523
rect 937 517 957 518
rect 937 514 957 515
rect 1253 526 1273 527
rect 1253 521 1273 522
rect 1691 525 1711 526
rect 1691 521 1707 525
rect 1965 522 1970 538
rect 1972 522 1978 542
rect 1980 526 1985 542
rect 1980 522 1981 526
rect 1993 538 1994 542
rect 1989 522 1994 538
rect 1996 522 2002 542
rect 2004 526 2009 542
rect 2004 522 2005 526
rect 2019 538 2020 542
rect 2015 522 2020 538
rect 2022 526 2027 542
rect 2022 522 2023 526
rect 2037 538 2038 542
rect 2033 522 2038 538
rect 2040 526 2045 542
rect 2040 522 2041 526
rect 2062 538 2063 542
rect 2058 522 2063 538
rect 2065 526 2070 542
rect 2065 522 2066 526
rect 2087 538 2088 542
rect 2083 522 2088 538
rect 2090 526 2095 542
rect 2090 522 2091 526
rect 1253 518 1273 519
rect 1253 513 1273 514
rect 1253 510 1273 511
rect -73 499 -72 503
rect 1691 501 1707 505
rect 1691 500 1711 501
rect 1691 497 1711 498
rect 1691 493 1693 497
rect 1697 493 1711 497
rect 1691 491 1711 493
rect 93 483 109 487
rect 1691 488 1711 489
rect 1695 484 1711 488
rect 93 482 113 483
rect 93 479 113 480
rect 97 475 113 479
rect 900 462 920 463
rect 900 459 920 460
rect 900 454 920 455
rect 900 451 920 452
rect 92 401 108 405
rect 88 400 108 401
rect 88 397 108 398
rect 88 393 104 397
rect 1969 391 1970 395
rect -200 375 -199 379
rect -204 359 -199 375
rect -197 359 -191 379
rect -189 363 -184 379
rect -189 359 -188 363
rect -176 375 -175 379
rect -180 359 -175 375
rect -173 359 -167 379
rect -165 363 -160 379
rect -165 359 -164 363
rect -150 375 -149 379
rect -154 359 -149 375
rect -147 363 -142 379
rect -147 359 -146 363
rect -132 375 -131 379
rect -136 359 -131 375
rect -129 363 -124 379
rect -129 359 -128 363
rect -107 375 -106 379
rect -111 359 -106 375
rect -104 363 -99 379
rect -104 359 -103 363
rect -82 375 -81 379
rect -86 359 -81 375
rect -79 363 -74 379
rect 1695 379 1711 383
rect 1691 378 1711 379
rect 88 373 104 377
rect 88 372 108 373
rect -79 359 -78 363
rect 88 369 108 370
rect 88 365 90 369
rect 94 365 108 369
rect 1691 375 1711 376
rect 1965 375 1970 391
rect 1972 375 1978 395
rect 1980 379 1985 395
rect 1980 375 1981 379
rect 1993 391 1994 395
rect 1989 375 1994 391
rect 1996 375 2002 395
rect 2004 379 2009 395
rect 2004 375 2005 379
rect 2019 391 2020 395
rect 2015 375 2020 391
rect 2022 379 2027 395
rect 2022 375 2023 379
rect 2037 391 2038 395
rect 2033 375 2038 391
rect 2040 379 2045 395
rect 2040 375 2041 379
rect 2062 391 2063 395
rect 2058 375 2063 391
rect 2065 379 2070 395
rect 2065 375 2066 379
rect 2087 391 2088 395
rect 2083 375 2088 391
rect 2090 379 2095 395
rect 2090 375 2091 379
rect 1691 371 1707 375
rect 938 370 958 371
rect 88 363 108 365
rect 88 360 108 361
rect 92 356 108 360
rect 938 367 958 368
rect 938 362 958 363
rect 938 359 958 360
rect 938 354 958 355
rect 1255 355 1275 356
rect 938 351 958 352
rect 1255 352 1275 353
rect 1691 351 1707 355
rect 1691 350 1711 351
rect 1255 347 1275 348
rect 1255 344 1275 345
rect 1255 339 1275 340
rect 1691 347 1711 348
rect 1691 343 1693 347
rect 1697 343 1711 347
rect 1691 341 1711 343
rect 1255 336 1275 337
rect 1691 338 1711 339
rect 1695 334 1711 338
rect 67 310 87 311
rect 67 307 87 308
rect 67 302 87 303
rect 67 299 87 300
rect -200 292 -199 296
rect -204 276 -199 292
rect -197 276 -191 296
rect -189 280 -184 296
rect -189 276 -188 280
rect -176 292 -175 296
rect -180 276 -175 292
rect -173 276 -167 296
rect -165 280 -160 296
rect -165 276 -164 280
rect -150 292 -149 296
rect -154 276 -149 292
rect -147 280 -142 296
rect -147 276 -146 280
rect -132 292 -131 296
rect -136 276 -131 292
rect -129 280 -124 296
rect -129 276 -128 280
rect -107 292 -106 296
rect -111 276 -106 292
rect -104 280 -99 296
rect -104 276 -103 280
rect -82 292 -81 296
rect -86 276 -81 292
rect -79 280 -74 296
rect 901 299 921 300
rect 901 296 921 297
rect 901 291 921 292
rect 901 288 921 289
rect -79 276 -78 280
rect 93 267 109 271
rect 93 266 113 267
rect 93 263 113 264
rect 97 259 113 263
rect 1695 241 1711 245
rect 1691 240 1711 241
rect 1970 244 1971 248
rect 1691 237 1711 238
rect 1691 233 1707 237
rect 1966 228 1971 244
rect 1973 228 1979 248
rect 1981 232 1986 248
rect 1981 228 1982 232
rect 1994 244 1995 248
rect 1990 228 1995 244
rect 1997 228 2003 248
rect 2005 232 2010 248
rect 2005 228 2006 232
rect 2020 244 2021 248
rect 2016 228 2021 244
rect 2023 232 2028 248
rect 2023 228 2024 232
rect 2038 244 2039 248
rect 2034 228 2039 244
rect 2041 232 2046 248
rect 2041 228 2042 232
rect 2063 244 2064 248
rect 2059 228 2064 244
rect 2066 232 2071 248
rect 2066 228 2067 232
rect 2088 244 2089 248
rect 2084 228 2089 244
rect 2091 232 2096 248
rect 2091 228 2092 232
rect 899 216 919 217
rect 899 213 919 214
rect 899 208 919 209
rect 1215 215 1235 216
rect 1215 212 1235 213
rect 899 205 919 206
rect 1215 207 1235 208
rect 1691 213 1707 217
rect 1691 212 1711 213
rect 1215 204 1235 205
rect 1691 209 1711 210
rect 1691 205 1693 209
rect 1697 205 1711 209
rect 1691 203 1711 205
rect 1691 200 1711 201
rect 1695 196 1711 200
rect 92 185 108 189
rect 88 184 108 185
rect 88 181 108 182
rect 88 177 104 181
rect -213 162 -212 166
rect -217 146 -212 162
rect -210 146 -204 166
rect -202 150 -197 166
rect -202 146 -201 150
rect -189 162 -188 166
rect -193 146 -188 162
rect -186 146 -180 166
rect -178 150 -173 166
rect -178 146 -177 150
rect -163 162 -162 166
rect -167 146 -162 162
rect -160 150 -155 166
rect -160 146 -159 150
rect -145 162 -144 166
rect -149 146 -144 162
rect -142 150 -137 166
rect -142 146 -141 150
rect -120 162 -119 166
rect -124 146 -119 162
rect -117 150 -112 166
rect -117 146 -116 150
rect -95 162 -94 166
rect -99 146 -94 162
rect -92 150 -87 166
rect 88 157 104 161
rect 88 156 108 157
rect -92 146 -91 150
rect 88 153 108 154
rect 88 149 90 153
rect 94 149 108 153
rect 88 147 108 149
rect 88 144 108 145
rect 92 140 108 144
rect 1970 139 1971 143
rect 1966 123 1971 139
rect 1973 123 1979 143
rect 1981 127 1986 143
rect 1981 123 1982 127
rect 1994 139 1995 143
rect 1990 123 1995 139
rect 1997 123 2003 143
rect 2005 127 2010 143
rect 2005 123 2006 127
rect 2020 139 2021 143
rect 2016 123 2021 139
rect 2023 127 2028 143
rect 2023 123 2024 127
rect 2038 139 2039 143
rect 2034 123 2039 139
rect 2041 127 2046 143
rect 2041 123 2042 127
rect 2063 139 2064 143
rect 2059 123 2064 139
rect 2066 127 2071 143
rect 2066 123 2067 127
rect 2088 139 2089 143
rect 2084 123 2089 139
rect 2091 127 2096 143
rect 2091 123 2092 127
rect 67 94 87 95
rect 67 91 87 92
rect 67 86 87 87
rect 67 83 87 84
rect -213 79 -212 83
rect -217 63 -212 79
rect -210 63 -204 83
rect -202 67 -197 83
rect -202 63 -201 67
rect -189 79 -188 83
rect -193 63 -188 79
rect -186 63 -180 83
rect -178 67 -173 83
rect -178 63 -177 67
rect -163 79 -162 83
rect -167 63 -162 79
rect -160 67 -155 83
rect -160 63 -159 67
rect -145 79 -144 83
rect -149 63 -144 79
rect -142 67 -137 83
rect -142 63 -141 67
rect -120 79 -119 83
rect -124 63 -119 79
rect -117 67 -112 83
rect -117 63 -116 67
rect -95 79 -94 83
rect -99 63 -94 79
rect -92 67 -87 83
rect -92 63 -91 67
rect 93 51 109 55
rect 93 50 113 51
rect 93 47 113 48
rect 97 43 113 47
<< ndcontact >>
rect 66 1049 70 1053
rect 66 1041 70 1045
rect 65 1021 69 1025
rect 71 1013 75 1017
rect -199 974 -195 978
rect -191 990 -187 994
rect -175 974 -171 978
rect -167 990 -163 994
rect -149 980 -145 984
rect -141 986 -137 990
rect -131 974 -127 978
rect -114 990 -110 994
rect -106 974 -102 978
rect -89 990 -85 994
rect 71 1004 75 1008
rect -81 980 -77 984
rect -73 986 -69 990
rect 900 979 950 983
rect 900 971 950 975
rect 900 963 950 967
rect 101 959 121 963
rect 900 955 950 959
rect 101 951 121 955
rect 900 947 950 951
rect 101 943 121 947
rect 900 939 950 943
rect -199 891 -195 895
rect -191 907 -187 911
rect -175 891 -171 895
rect -167 907 -163 911
rect -149 897 -145 901
rect -141 903 -137 907
rect -131 891 -127 895
rect -114 907 -110 911
rect -106 891 -102 895
rect -89 907 -85 911
rect 71 915 75 919
rect 77 907 81 911
rect -81 897 -77 901
rect -73 903 -69 907
rect 893 884 933 888
rect 893 876 933 880
rect 1969 874 1973 878
rect 1977 890 1981 894
rect 893 868 933 872
rect 1993 874 1997 878
rect 2001 890 2005 894
rect 893 860 933 864
rect 2019 880 2023 884
rect 2027 886 2031 890
rect 2037 874 2041 878
rect 2054 890 2058 894
rect 2062 874 2066 878
rect 2079 890 2083 894
rect 2087 880 2091 884
rect 2095 886 2099 890
rect 893 852 933 856
rect 1195 840 1245 844
rect 66 833 70 837
rect 1195 832 1245 836
rect 66 825 70 829
rect 1677 829 1681 833
rect 1195 824 1245 828
rect 1677 821 1681 825
rect 1195 816 1245 820
rect 65 805 69 809
rect 1195 808 1245 812
rect 71 797 75 801
rect 1195 800 1245 804
rect 1676 801 1680 805
rect -197 759 -193 763
rect -189 775 -185 779
rect -173 759 -169 763
rect -165 775 -161 779
rect -147 765 -143 769
rect -139 771 -135 775
rect -129 759 -125 763
rect -112 775 -108 779
rect -104 759 -100 763
rect -87 775 -83 779
rect 71 788 75 792
rect 888 789 918 793
rect 1682 793 1686 797
rect 888 781 918 785
rect 1682 784 1686 788
rect 1973 787 1977 791
rect 1981 803 1985 807
rect 1997 787 2001 791
rect 2005 803 2009 807
rect -79 765 -75 769
rect -71 771 -67 775
rect 888 773 918 777
rect 2023 793 2027 797
rect 2031 799 2035 803
rect 2041 787 2045 791
rect 2058 803 2062 807
rect 2066 787 2070 791
rect 2083 803 2087 807
rect 2091 793 2095 797
rect 2099 799 2103 803
rect 888 765 918 769
rect 101 743 121 747
rect 101 735 121 739
rect 101 727 121 731
rect 934 715 954 719
rect -197 676 -193 680
rect -189 692 -185 696
rect -173 676 -169 680
rect -165 692 -161 696
rect -147 682 -143 686
rect -139 688 -135 692
rect -129 676 -125 680
rect -112 692 -108 696
rect -104 676 -100 680
rect -87 692 -83 696
rect 934 707 954 711
rect 71 699 75 703
rect 934 699 954 703
rect -79 682 -75 686
rect -71 688 -67 692
rect 77 691 81 695
rect 66 617 70 621
rect 895 619 935 623
rect 66 609 70 613
rect 895 611 935 615
rect 895 603 935 607
rect 65 589 69 593
rect 895 595 935 599
rect 895 587 935 591
rect -198 550 -194 554
rect -190 566 -186 570
rect -174 550 -170 554
rect -166 566 -162 570
rect -148 556 -144 560
rect -140 562 -136 566
rect -130 550 -126 554
rect -113 566 -109 570
rect -105 550 -101 554
rect -88 566 -84 570
rect 71 581 75 585
rect 71 572 75 576
rect -80 556 -76 560
rect -72 562 -68 566
rect 1201 538 1241 542
rect 890 534 920 538
rect 101 527 121 531
rect 890 526 920 530
rect 101 519 121 523
rect 1201 530 1241 534
rect 1669 529 1673 533
rect 890 518 920 522
rect 101 511 121 515
rect 1201 522 1241 526
rect 890 510 920 514
rect 1669 521 1673 525
rect 1201 514 1241 518
rect 1201 506 1241 510
rect 1668 501 1672 505
rect -198 467 -194 471
rect -190 483 -186 487
rect -174 467 -170 471
rect -166 483 -162 487
rect -148 473 -144 477
rect -140 479 -136 483
rect -130 467 -126 471
rect -113 483 -109 487
rect -105 467 -101 471
rect -88 483 -84 487
rect 1674 493 1678 497
rect 1965 490 1969 494
rect 1973 506 1977 510
rect 71 483 75 487
rect -80 473 -76 477
rect -72 479 -68 483
rect 1674 484 1678 488
rect 1989 490 1993 494
rect 1997 506 2001 510
rect 77 475 81 479
rect 2015 496 2019 500
rect 2023 502 2027 506
rect 2033 490 2037 494
rect 2050 506 2054 510
rect 2058 490 2062 494
rect 2075 506 2079 510
rect 2083 496 2087 500
rect 2091 502 2095 506
rect 934 463 954 467
rect 934 455 954 459
rect 934 447 954 451
rect 66 401 70 405
rect 66 393 70 397
rect 1669 379 1673 383
rect 65 373 69 377
rect 891 371 921 375
rect 71 365 75 369
rect 1669 371 1673 375
rect 891 363 921 367
rect -204 327 -200 331
rect -196 343 -192 347
rect -180 327 -176 331
rect -172 343 -168 347
rect -154 333 -150 337
rect -146 339 -142 343
rect -136 327 -132 331
rect -119 343 -115 347
rect -111 327 -107 331
rect -94 343 -90 347
rect 71 356 75 360
rect 891 355 921 359
rect 1208 356 1238 360
rect 891 347 921 351
rect 1208 348 1238 352
rect 1668 351 1672 355
rect -86 333 -82 337
rect -78 339 -74 343
rect 1208 340 1238 344
rect 1674 343 1678 347
rect 1965 343 1969 347
rect 1973 359 1977 363
rect 1208 332 1238 336
rect 1674 334 1678 338
rect 1989 343 1993 347
rect 1997 359 2001 363
rect 2015 349 2019 353
rect 2023 355 2027 359
rect 2033 343 2037 347
rect 2050 359 2054 363
rect 2058 343 2062 347
rect 2075 359 2079 363
rect 2083 349 2087 353
rect 2091 355 2095 359
rect 101 311 121 315
rect 101 303 121 307
rect 101 295 121 299
rect 935 300 955 304
rect 935 292 955 296
rect 935 284 955 288
rect -204 244 -200 248
rect -196 260 -192 264
rect -180 244 -176 248
rect -172 260 -168 264
rect -154 250 -150 254
rect -146 256 -142 260
rect -136 244 -132 248
rect -119 260 -115 264
rect -111 244 -107 248
rect -94 260 -90 264
rect 71 267 75 271
rect -86 250 -82 254
rect -78 256 -74 260
rect 77 259 81 263
rect 1669 241 1673 245
rect 1669 233 1673 237
rect 933 217 953 221
rect 933 209 953 213
rect 1249 216 1269 220
rect 1668 213 1672 217
rect 933 201 953 205
rect 1249 208 1269 212
rect 1249 200 1269 204
rect 1674 205 1678 209
rect 1674 196 1678 200
rect 1966 196 1970 200
rect 1974 212 1978 216
rect 66 185 70 189
rect 1990 196 1994 200
rect 1998 212 2002 216
rect 2016 202 2020 206
rect 2024 208 2028 212
rect 2034 196 2038 200
rect 2051 212 2055 216
rect 2059 196 2063 200
rect 2076 212 2080 216
rect 2084 202 2088 206
rect 2092 208 2096 212
rect 66 177 70 181
rect 65 157 69 161
rect 71 149 75 153
rect -217 114 -213 118
rect -209 130 -205 134
rect -193 114 -189 118
rect -185 130 -181 134
rect -167 120 -163 124
rect -159 126 -155 130
rect -149 114 -145 118
rect -132 130 -128 134
rect -124 114 -120 118
rect -107 130 -103 134
rect 71 140 75 144
rect -99 120 -95 124
rect -91 126 -87 130
rect 101 95 121 99
rect 1966 91 1970 95
rect 1974 107 1978 111
rect 101 87 121 91
rect 101 79 121 83
rect 1990 91 1994 95
rect 1998 107 2002 111
rect 2016 97 2020 101
rect 2024 103 2028 107
rect 2034 91 2038 95
rect 2051 107 2055 111
rect 2059 91 2063 95
rect 2076 107 2080 111
rect 2084 97 2088 101
rect 2092 103 2096 107
rect -217 31 -213 35
rect -209 47 -205 51
rect -193 31 -189 35
rect -185 47 -181 51
rect -167 37 -163 41
rect -159 43 -155 47
rect -149 31 -145 35
rect -132 47 -128 51
rect -124 31 -120 35
rect -107 47 -103 51
rect 71 51 75 55
rect -99 37 -95 41
rect -91 43 -87 47
rect 77 43 81 47
<< pdcontact >>
rect 88 1049 92 1053
rect 104 1041 108 1045
rect -199 1022 -195 1026
rect -183 1006 -179 1010
rect -175 1022 -171 1026
rect -159 1006 -155 1010
rect -149 1022 -145 1026
rect -141 1006 -137 1010
rect -131 1022 -127 1026
rect -123 1006 -119 1010
rect -106 1022 -102 1026
rect -98 1006 -94 1010
rect -81 1022 -77 1026
rect 104 1021 108 1025
rect -73 1006 -69 1010
rect 90 1013 94 1017
rect 88 1004 92 1008
rect 964 979 984 983
rect 964 971 984 975
rect 67 959 87 963
rect 964 963 984 967
rect 67 951 87 955
rect 964 955 984 959
rect 67 943 87 947
rect 964 947 984 951
rect -199 939 -195 943
rect -183 923 -179 927
rect -175 939 -171 943
rect -159 923 -155 927
rect -149 939 -145 943
rect -141 923 -137 927
rect -131 939 -127 943
rect -123 923 -119 927
rect -106 939 -102 943
rect -98 923 -94 927
rect -81 939 -77 943
rect 964 939 984 943
rect -73 923 -69 927
rect 1969 922 1973 926
rect 109 915 113 919
rect 93 907 97 911
rect 1985 906 1989 910
rect 1993 922 1997 926
rect 2009 906 2013 910
rect 2019 922 2023 926
rect 2027 906 2031 910
rect 2037 922 2041 926
rect 2045 906 2049 910
rect 2062 922 2066 926
rect 2070 906 2074 910
rect 2087 922 2091 926
rect 2095 906 2099 910
rect 945 884 965 888
rect 945 876 965 880
rect 945 868 965 872
rect 945 860 965 864
rect 945 852 965 856
rect 88 833 92 837
rect 1259 840 1279 844
rect 104 825 108 829
rect 1259 832 1279 836
rect 1973 835 1977 839
rect 1699 829 1703 833
rect 1259 824 1279 828
rect 1715 821 1719 825
rect 1259 816 1279 820
rect 1989 819 1993 823
rect 1997 835 2001 839
rect 2013 819 2017 823
rect 2023 835 2027 839
rect 2031 819 2035 823
rect 2041 835 2045 839
rect 2049 819 2053 823
rect 2066 835 2070 839
rect 2074 819 2078 823
rect 2091 835 2095 839
rect 2099 819 2103 823
rect -197 807 -193 811
rect -181 791 -177 795
rect -173 807 -169 811
rect -157 791 -153 795
rect -147 807 -143 811
rect -139 791 -135 795
rect -129 807 -125 811
rect -121 791 -117 795
rect -104 807 -100 811
rect -96 791 -92 795
rect -79 807 -75 811
rect 104 805 108 809
rect 1259 808 1279 812
rect -71 791 -67 795
rect 90 797 94 801
rect 1259 800 1279 804
rect 1715 801 1719 805
rect 88 788 92 792
rect 935 789 955 793
rect 1701 793 1705 797
rect 935 781 955 785
rect 1699 784 1703 788
rect 935 773 955 777
rect 935 765 955 769
rect 67 743 87 747
rect 67 735 87 739
rect -197 724 -193 728
rect -181 708 -177 712
rect -173 724 -169 728
rect -157 708 -153 712
rect -147 724 -143 728
rect -139 708 -135 712
rect -129 724 -125 728
rect -121 708 -117 712
rect -104 724 -100 728
rect -96 708 -92 712
rect -79 724 -75 728
rect 67 727 87 731
rect 900 715 920 719
rect -71 708 -67 712
rect 900 707 920 711
rect 109 699 113 703
rect 900 699 920 703
rect 93 691 97 695
rect 88 617 92 621
rect 947 619 967 623
rect 104 609 108 613
rect 947 611 967 615
rect -198 598 -194 602
rect -182 582 -178 586
rect -174 598 -170 602
rect -158 582 -154 586
rect -148 598 -144 602
rect -140 582 -136 586
rect -130 598 -126 602
rect -122 582 -118 586
rect -105 598 -101 602
rect -97 582 -93 586
rect -80 598 -76 602
rect 947 603 967 607
rect 104 589 108 593
rect 947 595 967 599
rect 947 587 967 591
rect -72 582 -68 586
rect 90 581 94 585
rect 88 572 92 576
rect 67 527 87 531
rect 937 534 957 538
rect 1253 538 1273 542
rect 1965 538 1969 542
rect 67 519 87 523
rect -198 515 -194 519
rect -182 499 -178 503
rect -174 515 -170 519
rect -158 499 -154 503
rect -148 515 -144 519
rect -140 499 -136 503
rect -130 515 -126 519
rect -122 499 -118 503
rect -105 515 -101 519
rect -97 499 -93 503
rect -80 515 -76 519
rect 937 526 957 530
rect 1253 530 1273 534
rect 1691 529 1695 533
rect 67 511 87 515
rect 937 518 957 522
rect 1253 522 1273 526
rect 1707 521 1711 525
rect 1981 522 1985 526
rect 1989 538 1993 542
rect 2005 522 2009 526
rect 2015 538 2019 542
rect 2023 522 2027 526
rect 2033 538 2037 542
rect 2041 522 2045 526
rect 2058 538 2062 542
rect 2066 522 2070 526
rect 2083 538 2087 542
rect 2091 522 2095 526
rect 937 510 957 514
rect 1253 514 1273 518
rect 1253 506 1273 510
rect -72 499 -68 503
rect 1707 501 1711 505
rect 1693 493 1697 497
rect 109 483 113 487
rect 1691 484 1695 488
rect 93 475 97 479
rect 900 463 920 467
rect 900 455 920 459
rect 900 447 920 451
rect 88 401 92 405
rect 104 393 108 397
rect 1965 391 1969 395
rect -204 375 -200 379
rect -188 359 -184 363
rect -180 375 -176 379
rect -164 359 -160 363
rect -154 375 -150 379
rect -146 359 -142 363
rect -136 375 -132 379
rect -128 359 -124 363
rect -111 375 -107 379
rect -103 359 -99 363
rect -86 375 -82 379
rect 1691 379 1695 383
rect 104 373 108 377
rect -78 359 -74 363
rect 90 365 94 369
rect 938 371 958 375
rect 1981 375 1985 379
rect 1989 391 1993 395
rect 2005 375 2009 379
rect 2015 391 2019 395
rect 2023 375 2027 379
rect 2033 391 2037 395
rect 2041 375 2045 379
rect 2058 391 2062 395
rect 2066 375 2070 379
rect 2083 391 2087 395
rect 2091 375 2095 379
rect 1707 371 1711 375
rect 88 356 92 360
rect 938 363 958 367
rect 938 355 958 359
rect 1255 356 1275 360
rect 938 347 958 351
rect 1255 348 1275 352
rect 1707 351 1711 355
rect 1255 340 1275 344
rect 1693 343 1697 347
rect 1255 332 1275 336
rect 1691 334 1695 338
rect 67 311 87 315
rect 67 303 87 307
rect 901 300 921 304
rect -204 292 -200 296
rect -188 276 -184 280
rect -180 292 -176 296
rect -164 276 -160 280
rect -154 292 -150 296
rect -146 276 -142 280
rect -136 292 -132 296
rect -128 276 -124 280
rect -111 292 -107 296
rect -103 276 -99 280
rect -86 292 -82 296
rect 67 295 87 299
rect 901 292 921 296
rect 901 284 921 288
rect -78 276 -74 280
rect 109 267 113 271
rect 93 259 97 263
rect 1691 241 1695 245
rect 1966 244 1970 248
rect 1707 233 1711 237
rect 1982 228 1986 232
rect 1990 244 1994 248
rect 2006 228 2010 232
rect 2016 244 2020 248
rect 2024 228 2028 232
rect 2034 244 2038 248
rect 2042 228 2046 232
rect 2059 244 2063 248
rect 2067 228 2071 232
rect 2084 244 2088 248
rect 2092 228 2096 232
rect 899 217 919 221
rect 1215 216 1235 220
rect 899 209 919 213
rect 1215 208 1235 212
rect 899 201 919 205
rect 1707 213 1711 217
rect 1215 200 1235 204
rect 1693 205 1697 209
rect 1691 196 1695 200
rect 88 185 92 189
rect 104 177 108 181
rect -217 162 -213 166
rect -201 146 -197 150
rect -193 162 -189 166
rect -177 146 -173 150
rect -167 162 -163 166
rect -159 146 -155 150
rect -149 162 -145 166
rect -141 146 -137 150
rect -124 162 -120 166
rect -116 146 -112 150
rect -99 162 -95 166
rect 104 157 108 161
rect -91 146 -87 150
rect 90 149 94 153
rect 88 140 92 144
rect 1966 139 1970 143
rect 1982 123 1986 127
rect 1990 139 1994 143
rect 2006 123 2010 127
rect 2016 139 2020 143
rect 2024 123 2028 127
rect 2034 139 2038 143
rect 2042 123 2046 127
rect 2059 139 2063 143
rect 2067 123 2071 127
rect 2084 139 2088 143
rect 2092 123 2096 127
rect 67 95 87 99
rect 67 87 87 91
rect -217 79 -213 83
rect -201 63 -197 67
rect -193 79 -189 83
rect -177 63 -173 67
rect -167 79 -163 83
rect -159 63 -155 67
rect -149 79 -145 83
rect -141 63 -137 67
rect -124 79 -120 83
rect -116 63 -112 67
rect -99 79 -95 83
rect 67 79 87 83
rect -91 63 -87 67
rect 109 51 113 55
rect 93 43 97 47
<< polysilicon >>
rect 62 1046 66 1048
rect 76 1046 88 1048
rect 108 1046 112 1048
rect -194 1026 -192 1030
rect -186 1026 -184 1030
rect -170 1026 -168 1030
rect -162 1026 -160 1030
rect -144 1026 -142 1030
rect -126 1026 -124 1029
rect -101 1026 -99 1029
rect -76 1026 -74 1030
rect 62 1018 65 1020
rect 75 1018 88 1020
rect 108 1018 111 1020
rect 58 1010 59 1011
rect 63 1010 65 1011
rect 58 1009 65 1010
rect 75 1009 79 1011
rect 82 1009 88 1011
rect 108 1009 120 1011
rect -194 994 -192 1006
rect -194 971 -192 974
rect -186 965 -184 1006
rect -170 994 -168 1006
rect -170 971 -168 974
rect -185 962 -184 965
rect -162 962 -160 1006
rect -144 990 -142 1006
rect -126 994 -124 1006
rect -117 994 -115 998
rect -101 994 -99 1006
rect -92 994 -90 998
rect -144 976 -142 980
rect -76 990 -74 1006
rect -76 976 -74 980
rect 892 976 900 978
rect 950 976 964 978
rect 984 976 987 978
rect -126 969 -124 974
rect -117 961 -115 974
rect -101 969 -99 974
rect -92 961 -90 974
rect 892 968 900 970
rect 950 968 964 970
rect 984 968 987 970
rect 892 960 900 962
rect 950 960 964 962
rect 984 960 987 962
rect 54 956 67 958
rect 87 956 101 958
rect 121 956 126 958
rect 892 952 900 954
rect 950 952 964 954
rect 984 952 987 954
rect 54 948 67 950
rect 87 948 101 950
rect 121 948 126 950
rect -194 943 -192 947
rect -186 943 -184 947
rect -170 943 -168 947
rect -162 943 -160 947
rect -144 943 -142 947
rect -126 943 -124 946
rect -101 943 -99 946
rect -76 943 -74 947
rect 892 944 900 946
rect 950 944 964 946
rect 984 944 987 946
rect 1974 926 1976 930
rect 1982 926 1984 930
rect 1998 926 2000 930
rect 2006 926 2008 930
rect 2024 926 2026 930
rect 2042 926 2044 929
rect 2067 926 2069 929
rect 2092 926 2094 930
rect -194 911 -192 923
rect -194 888 -192 891
rect -186 882 -184 923
rect -170 911 -168 923
rect -170 888 -168 891
rect -185 879 -184 882
rect -162 879 -160 923
rect -144 907 -142 923
rect -126 911 -124 923
rect -117 911 -115 915
rect -101 911 -99 923
rect -92 911 -90 915
rect -144 893 -142 897
rect -76 907 -74 923
rect 67 912 71 914
rect 81 912 93 914
rect 113 912 117 914
rect -76 893 -74 897
rect 1974 894 1976 906
rect -126 886 -124 891
rect -117 877 -115 891
rect -101 886 -99 891
rect -92 877 -90 891
rect 888 881 893 883
rect 933 881 945 883
rect 965 881 968 883
rect 888 873 893 875
rect 933 873 945 875
rect 965 873 968 875
rect 1974 871 1976 874
rect 888 865 893 867
rect 933 865 945 867
rect 965 865 968 867
rect 1982 865 1984 906
rect 1998 894 2000 906
rect 1998 871 2000 874
rect 1983 862 1984 865
rect 2006 862 2008 906
rect 2024 890 2026 906
rect 2042 894 2044 906
rect 2051 894 2053 898
rect 2067 894 2069 906
rect 2076 894 2078 898
rect 2024 876 2026 880
rect 2092 890 2094 906
rect 2092 876 2094 880
rect 2042 869 2044 874
rect 2051 860 2053 874
rect 2067 869 2069 874
rect 2076 860 2078 874
rect 888 857 893 859
rect 933 857 945 859
rect 965 857 968 859
rect 1978 839 1980 843
rect 1986 839 1988 843
rect 2002 839 2004 843
rect 2010 839 2012 843
rect 2028 839 2030 843
rect 2046 839 2048 842
rect 2071 839 2073 842
rect 2096 839 2098 843
rect 1187 837 1195 839
rect 1245 837 1259 839
rect 1279 837 1282 839
rect 62 830 66 832
rect 76 830 88 832
rect 108 830 112 832
rect 1187 829 1195 831
rect 1245 829 1259 831
rect 1279 829 1282 831
rect 1673 826 1677 828
rect 1687 826 1699 828
rect 1719 826 1723 828
rect 1187 821 1195 823
rect 1245 821 1259 823
rect 1279 821 1282 823
rect -192 811 -190 815
rect -184 811 -182 815
rect -168 811 -166 815
rect -160 811 -158 815
rect -142 811 -140 815
rect -124 811 -122 814
rect -99 811 -97 814
rect -74 811 -72 815
rect 1187 813 1195 815
rect 1245 813 1259 815
rect 1279 813 1282 815
rect 1978 807 1980 819
rect 1187 805 1195 807
rect 1245 805 1259 807
rect 1279 805 1282 807
rect 62 802 65 804
rect 75 802 88 804
rect 108 802 111 804
rect 58 794 59 795
rect 1673 798 1676 800
rect 1686 798 1699 800
rect 1719 798 1722 800
rect 63 794 65 795
rect 58 793 65 794
rect 75 793 79 795
rect 82 793 88 795
rect 108 793 120 795
rect -192 779 -190 791
rect -192 756 -190 759
rect -184 750 -182 791
rect -168 779 -166 791
rect -168 756 -166 759
rect -183 747 -182 750
rect -160 747 -158 791
rect -142 775 -140 791
rect -124 779 -122 791
rect -115 779 -113 783
rect -99 779 -97 791
rect -90 779 -88 783
rect -142 761 -140 765
rect -74 775 -72 791
rect 1669 790 1670 791
rect 1674 790 1676 791
rect 1669 789 1676 790
rect 1686 789 1690 791
rect 1693 789 1699 791
rect 1719 789 1731 791
rect 885 786 888 788
rect 918 786 935 788
rect 955 786 958 788
rect 1978 784 1980 787
rect 885 778 888 780
rect 918 778 935 780
rect 955 778 958 780
rect 1986 778 1988 819
rect 2002 807 2004 819
rect 2002 784 2004 787
rect 1987 775 1988 778
rect 2010 775 2012 819
rect 2028 803 2030 819
rect 2046 807 2048 819
rect 2055 807 2057 811
rect 2071 807 2073 819
rect 2080 807 2082 811
rect 2028 789 2030 793
rect 2096 803 2098 819
rect 2096 789 2098 793
rect 2046 782 2048 787
rect 2055 773 2057 787
rect 2071 782 2073 787
rect 2080 773 2082 787
rect 885 770 888 772
rect 918 770 935 772
rect 955 770 958 772
rect -74 761 -72 765
rect -124 754 -122 759
rect -115 746 -113 759
rect -99 754 -97 759
rect -90 746 -88 759
rect 54 740 67 742
rect 87 740 101 742
rect 121 740 126 742
rect -192 728 -190 732
rect -184 728 -182 732
rect -168 728 -166 732
rect -160 728 -158 732
rect -142 728 -140 732
rect -124 728 -122 731
rect -99 728 -97 731
rect -74 728 -72 732
rect 54 732 67 734
rect 87 732 101 734
rect 121 732 126 734
rect 887 712 900 714
rect 920 712 934 714
rect 954 712 959 714
rect -192 696 -190 708
rect -192 673 -190 676
rect -184 667 -182 708
rect -168 696 -166 708
rect -168 673 -166 676
rect -183 664 -182 667
rect -160 664 -158 708
rect -142 692 -140 708
rect -124 696 -122 708
rect -115 696 -113 700
rect -99 696 -97 708
rect -90 696 -88 700
rect -142 678 -140 682
rect -74 692 -72 708
rect 887 704 900 706
rect 920 704 934 706
rect 954 704 959 706
rect 67 696 71 698
rect 81 696 93 698
rect 113 696 117 698
rect -74 678 -72 682
rect -124 671 -122 676
rect -115 662 -113 676
rect -99 671 -97 676
rect -90 662 -88 676
rect 62 614 66 616
rect 76 614 88 616
rect 108 614 112 616
rect 890 616 895 618
rect 935 616 947 618
rect 967 616 970 618
rect 890 608 895 610
rect 935 608 947 610
rect 967 608 970 610
rect -193 602 -191 606
rect -185 602 -183 606
rect -169 602 -167 606
rect -161 602 -159 606
rect -143 602 -141 606
rect -125 602 -123 605
rect -100 602 -98 605
rect -75 602 -73 606
rect 890 600 895 602
rect 935 600 947 602
rect 967 600 970 602
rect 890 592 895 594
rect 935 592 947 594
rect 967 592 970 594
rect 62 586 65 588
rect 75 586 88 588
rect 108 586 111 588
rect -193 570 -191 582
rect -193 547 -191 550
rect -185 541 -183 582
rect -169 570 -167 582
rect -169 547 -167 550
rect -184 538 -183 541
rect -161 538 -159 582
rect -143 566 -141 582
rect -125 570 -123 582
rect -116 570 -114 574
rect -100 570 -98 582
rect -91 570 -89 574
rect -143 552 -141 556
rect -75 566 -73 582
rect 58 578 59 579
rect 63 578 65 579
rect 58 577 65 578
rect 75 577 79 579
rect 82 577 88 579
rect 108 577 120 579
rect -75 552 -73 556
rect -125 545 -123 550
rect -116 537 -114 550
rect -100 545 -98 550
rect -91 537 -89 550
rect 1970 542 1972 546
rect 1978 542 1980 546
rect 1994 542 1996 546
rect 2002 542 2004 546
rect 2020 542 2022 546
rect 2038 542 2040 545
rect 2063 542 2065 545
rect 2088 542 2090 546
rect 1196 535 1201 537
rect 1241 535 1253 537
rect 1273 535 1276 537
rect 887 531 890 533
rect 920 531 937 533
rect 957 531 960 533
rect 54 524 67 526
rect 87 524 101 526
rect 121 524 126 526
rect -193 519 -191 523
rect -185 519 -183 523
rect -169 519 -167 523
rect -161 519 -159 523
rect -143 519 -141 523
rect -125 519 -123 522
rect -100 519 -98 522
rect -75 519 -73 523
rect 1196 527 1201 529
rect 1241 527 1253 529
rect 1273 527 1276 529
rect 887 523 890 525
rect 920 523 937 525
rect 957 523 960 525
rect 54 516 67 518
rect 87 516 101 518
rect 121 516 126 518
rect 887 515 890 517
rect 920 515 937 517
rect 957 515 960 517
rect 1665 526 1669 528
rect 1679 526 1691 528
rect 1711 526 1715 528
rect 1196 519 1201 521
rect 1241 519 1253 521
rect 1273 519 1276 521
rect 1196 511 1201 513
rect 1241 511 1253 513
rect 1273 511 1276 513
rect 1970 510 1972 522
rect -193 487 -191 499
rect -193 464 -191 467
rect -185 458 -183 499
rect -169 487 -167 499
rect -169 464 -167 467
rect -184 455 -183 458
rect -161 455 -159 499
rect -143 483 -141 499
rect -125 487 -123 499
rect -116 487 -114 491
rect -100 487 -98 499
rect -91 487 -89 491
rect -143 469 -141 473
rect -75 483 -73 499
rect 1665 498 1668 500
rect 1678 498 1691 500
rect 1711 498 1714 500
rect 1661 490 1662 491
rect 1666 490 1668 491
rect 1661 489 1668 490
rect 1678 489 1682 491
rect 1685 489 1691 491
rect 1711 489 1723 491
rect 1970 487 1972 490
rect 67 480 71 482
rect 81 480 93 482
rect 113 480 117 482
rect 1978 481 1980 522
rect 1994 510 1996 522
rect 1994 487 1996 490
rect 1979 478 1980 481
rect 2002 478 2004 522
rect 2020 506 2022 522
rect 2038 510 2040 522
rect 2047 510 2049 514
rect 2063 510 2065 522
rect 2072 510 2074 514
rect 2020 492 2022 496
rect 2088 506 2090 522
rect 2088 492 2090 496
rect 2038 485 2040 490
rect 2047 476 2049 490
rect 2063 485 2065 490
rect 2072 476 2074 490
rect -75 469 -73 473
rect -125 462 -123 467
rect -116 453 -114 467
rect -100 462 -98 467
rect -91 453 -89 467
rect 887 460 900 462
rect 920 460 934 462
rect 954 460 959 462
rect 887 452 900 454
rect 920 452 934 454
rect 954 452 959 454
rect 62 398 66 400
rect 76 398 88 400
rect 108 398 112 400
rect 1970 395 1972 399
rect 1978 395 1980 399
rect 1994 395 1996 399
rect 2002 395 2004 399
rect 2020 395 2022 399
rect 2038 395 2040 398
rect 2063 395 2065 398
rect 2088 395 2090 399
rect -199 379 -197 383
rect -191 379 -189 383
rect -175 379 -173 383
rect -167 379 -165 383
rect -149 379 -147 383
rect -131 379 -129 382
rect -106 379 -104 382
rect -81 379 -79 383
rect 1665 376 1669 378
rect 1679 376 1691 378
rect 1711 376 1715 378
rect 62 370 65 372
rect 75 370 88 372
rect 108 370 111 372
rect 58 362 59 363
rect 888 368 891 370
rect 921 368 938 370
rect 958 368 961 370
rect 63 362 65 363
rect 58 361 65 362
rect 75 361 79 363
rect 82 361 88 363
rect 108 361 120 363
rect -199 347 -197 359
rect -199 324 -197 327
rect -191 318 -189 359
rect -175 347 -173 359
rect -175 324 -173 327
rect -190 315 -189 318
rect -167 315 -165 359
rect -149 343 -147 359
rect -131 347 -129 359
rect -122 347 -120 351
rect -106 347 -104 359
rect -97 347 -95 351
rect -149 329 -147 333
rect -81 343 -79 359
rect 1970 363 1972 375
rect 888 360 891 362
rect 921 360 938 362
rect 958 360 961 362
rect 888 352 891 354
rect 921 352 938 354
rect 958 352 961 354
rect 1205 353 1208 355
rect 1238 353 1255 355
rect 1275 353 1278 355
rect 1665 348 1668 350
rect 1678 348 1691 350
rect 1711 348 1714 350
rect 1205 345 1208 347
rect 1238 345 1255 347
rect 1275 345 1278 347
rect 1661 340 1662 341
rect 1666 340 1668 341
rect 1661 339 1668 340
rect 1678 339 1682 341
rect 1685 339 1691 341
rect 1711 339 1723 341
rect 1970 340 1972 343
rect 1205 337 1208 339
rect 1238 337 1255 339
rect 1275 337 1278 339
rect -81 329 -79 333
rect 1978 334 1980 375
rect 1994 363 1996 375
rect 1994 340 1996 343
rect 1979 331 1980 334
rect 2002 331 2004 375
rect 2020 359 2022 375
rect 2038 363 2040 375
rect 2047 363 2049 367
rect 2063 363 2065 375
rect 2072 363 2074 367
rect 2020 345 2022 349
rect 2088 359 2090 375
rect 2088 345 2090 349
rect 2038 338 2040 343
rect 2047 329 2049 343
rect 2063 338 2065 343
rect 2072 329 2074 343
rect -131 322 -129 327
rect -122 314 -120 327
rect -106 322 -104 327
rect -97 314 -95 327
rect 54 308 67 310
rect 87 308 101 310
rect 121 308 126 310
rect -199 296 -197 300
rect -191 296 -189 300
rect -175 296 -173 300
rect -167 296 -165 300
rect -149 296 -147 300
rect -131 296 -129 299
rect -106 296 -104 299
rect -81 296 -79 300
rect 54 300 67 302
rect 87 300 101 302
rect 121 300 126 302
rect 888 297 901 299
rect 921 297 935 299
rect 955 297 960 299
rect 888 289 901 291
rect 921 289 935 291
rect 955 289 960 291
rect -199 264 -197 276
rect -199 241 -197 244
rect -191 235 -189 276
rect -175 264 -173 276
rect -175 241 -173 244
rect -190 232 -189 235
rect -167 232 -165 276
rect -149 260 -147 276
rect -131 264 -129 276
rect -122 264 -120 268
rect -106 264 -104 276
rect -97 264 -95 268
rect -149 246 -147 250
rect -81 260 -79 276
rect 67 264 71 266
rect 81 264 93 266
rect 113 264 117 266
rect -81 246 -79 250
rect 1971 248 1973 252
rect 1979 248 1981 252
rect 1995 248 1997 252
rect 2003 248 2005 252
rect 2021 248 2023 252
rect 2039 248 2041 251
rect 2064 248 2066 251
rect 2089 248 2091 252
rect -131 239 -129 244
rect -122 230 -120 244
rect -106 239 -104 244
rect -97 230 -95 244
rect 1665 238 1669 240
rect 1679 238 1691 240
rect 1711 238 1715 240
rect 886 214 899 216
rect 919 214 933 216
rect 953 214 958 216
rect 1202 213 1215 215
rect 1235 213 1249 215
rect 1269 213 1274 215
rect 886 206 899 208
rect 919 206 933 208
rect 953 206 958 208
rect 1971 216 1973 228
rect 1665 210 1668 212
rect 1678 210 1691 212
rect 1711 210 1714 212
rect 1202 205 1215 207
rect 1235 205 1249 207
rect 1269 205 1274 207
rect 1661 202 1662 203
rect 1666 202 1668 203
rect 1661 201 1668 202
rect 1678 201 1682 203
rect 1685 201 1691 203
rect 1711 201 1723 203
rect 1971 193 1973 196
rect 1979 187 1981 228
rect 1995 216 1997 228
rect 1995 193 1997 196
rect 62 182 66 184
rect 76 182 88 184
rect 108 182 112 184
rect 1980 184 1981 187
rect 2003 184 2005 228
rect 2021 212 2023 228
rect 2039 216 2041 228
rect 2048 216 2050 220
rect 2064 216 2066 228
rect 2073 216 2075 220
rect 2021 198 2023 202
rect 2089 212 2091 228
rect 2089 198 2091 202
rect 2039 191 2041 196
rect 2048 182 2050 196
rect 2064 191 2066 196
rect 2073 182 2075 196
rect -212 166 -210 170
rect -204 166 -202 170
rect -188 166 -186 170
rect -180 166 -178 170
rect -162 166 -160 170
rect -144 166 -142 169
rect -119 166 -117 169
rect -94 166 -92 170
rect 62 154 65 156
rect 75 154 88 156
rect 108 154 111 156
rect 58 146 59 147
rect 63 146 65 147
rect -212 134 -210 146
rect -212 111 -210 114
rect -204 105 -202 146
rect -188 134 -186 146
rect -188 111 -186 114
rect -203 102 -202 105
rect -180 102 -178 146
rect -162 130 -160 146
rect -144 134 -142 146
rect -135 134 -133 138
rect -119 134 -117 146
rect -110 134 -108 138
rect -162 116 -160 120
rect -94 130 -92 146
rect 58 145 65 146
rect 75 145 79 147
rect 82 145 88 147
rect 108 145 120 147
rect 1971 143 1973 147
rect 1979 143 1981 147
rect 1995 143 1997 147
rect 2003 143 2005 147
rect 2021 143 2023 147
rect 2039 143 2041 146
rect 2064 143 2066 146
rect 2089 143 2091 147
rect -94 116 -92 120
rect -144 109 -142 114
rect -135 101 -133 114
rect -119 109 -117 114
rect -110 101 -108 114
rect 1971 111 1973 123
rect 54 92 67 94
rect 87 92 101 94
rect 121 92 126 94
rect -212 83 -210 87
rect -204 83 -202 87
rect -188 83 -186 87
rect -180 83 -178 87
rect -162 83 -160 87
rect -144 83 -142 86
rect -119 83 -117 86
rect -94 83 -92 87
rect 1971 88 1973 91
rect 54 84 67 86
rect 87 84 101 86
rect 121 84 126 86
rect 1979 82 1981 123
rect 1995 111 1997 123
rect 1995 88 1997 91
rect 1980 79 1981 82
rect 2003 79 2005 123
rect 2021 107 2023 123
rect 2039 111 2041 123
rect 2048 111 2050 115
rect 2064 111 2066 123
rect 2073 111 2075 115
rect 2021 93 2023 97
rect 2089 107 2091 123
rect 2089 93 2091 97
rect 2039 86 2041 91
rect 2048 77 2050 91
rect 2064 86 2066 91
rect 2073 77 2075 91
rect -212 51 -210 63
rect -212 28 -210 31
rect -204 22 -202 63
rect -188 51 -186 63
rect -188 28 -186 31
rect -203 19 -202 22
rect -180 19 -178 63
rect -162 47 -160 63
rect -144 51 -142 63
rect -135 51 -133 55
rect -119 51 -117 63
rect -110 51 -108 55
rect -162 33 -160 37
rect -94 47 -92 63
rect 67 48 71 50
rect 81 48 93 50
rect 113 48 117 50
rect -94 33 -92 37
rect -144 26 -142 31
rect -135 17 -133 31
rect -119 26 -117 31
rect -110 17 -108 31
<< polycontact >>
rect 77 1042 81 1046
rect 77 1020 81 1024
rect 59 1010 63 1014
rect 115 1011 119 1015
rect -198 995 -194 999
rect -174 995 -170 999
rect -189 961 -185 965
rect -166 961 -162 965
rect -148 994 -144 998
rect -130 995 -126 999
rect -105 995 -101 999
rect -80 994 -76 998
rect 888 975 892 979
rect -121 961 -117 965
rect -96 961 -92 965
rect 888 967 892 971
rect 50 955 54 959
rect 888 959 892 963
rect 50 947 54 951
rect 888 951 892 955
rect 888 943 892 947
rect -198 912 -194 916
rect -174 912 -170 916
rect -189 878 -185 882
rect -166 878 -162 882
rect -148 911 -144 915
rect -130 912 -126 916
rect -105 912 -101 916
rect -80 911 -76 915
rect 82 914 86 918
rect 1970 895 1974 899
rect -121 878 -117 882
rect -96 878 -92 882
rect 884 880 888 884
rect 884 872 888 876
rect 884 864 888 868
rect 1994 895 1998 899
rect 884 856 888 860
rect 1979 861 1983 865
rect 2002 861 2006 865
rect 2020 894 2024 898
rect 2038 895 2042 899
rect 2063 895 2067 899
rect 2088 894 2092 898
rect 2047 861 2051 865
rect 2072 861 2076 865
rect 1183 836 1187 840
rect 77 826 81 830
rect 1183 828 1187 832
rect 1183 820 1187 824
rect 1688 822 1692 826
rect 1183 812 1187 816
rect 77 804 81 808
rect 1183 804 1187 808
rect 1974 808 1978 812
rect 59 794 63 798
rect 1688 800 1692 804
rect 115 795 119 799
rect -196 780 -192 784
rect -172 780 -168 784
rect -187 746 -183 750
rect -164 746 -160 750
rect -146 779 -142 783
rect -128 780 -124 784
rect -103 780 -99 784
rect -78 779 -74 783
rect 881 785 885 789
rect 1670 790 1674 794
rect 1726 791 1730 795
rect 881 777 885 781
rect 1998 808 2002 812
rect 881 769 885 773
rect 1983 774 1987 778
rect 2006 774 2010 778
rect 2024 807 2028 811
rect 2042 808 2046 812
rect 2067 808 2071 812
rect 2092 807 2096 811
rect 2051 774 2055 778
rect 2076 774 2080 778
rect -119 746 -115 750
rect -94 746 -90 750
rect 50 739 54 743
rect 50 731 54 735
rect 883 711 887 715
rect -196 697 -192 701
rect -172 697 -168 701
rect -187 663 -183 667
rect -164 663 -160 667
rect -146 696 -142 700
rect -128 697 -124 701
rect -103 697 -99 701
rect -78 696 -74 700
rect 883 703 887 707
rect 82 698 86 702
rect -119 663 -115 667
rect -94 663 -90 667
rect 886 615 890 619
rect 77 610 81 614
rect 886 607 890 611
rect 886 599 890 603
rect 77 588 81 592
rect 886 591 890 595
rect -197 571 -193 575
rect -173 571 -169 575
rect -188 537 -184 541
rect -165 537 -161 541
rect -147 570 -143 574
rect -129 571 -125 575
rect -104 571 -100 575
rect -79 570 -75 574
rect 59 578 63 582
rect 115 579 119 583
rect -120 537 -116 541
rect -95 537 -91 541
rect 50 523 54 527
rect 883 530 887 534
rect 1192 534 1196 538
rect 50 515 54 519
rect 883 522 887 526
rect 1192 526 1196 530
rect 883 514 887 518
rect 1192 518 1196 522
rect 1680 522 1684 526
rect 1192 510 1196 514
rect 1966 511 1970 515
rect 1680 500 1684 504
rect -197 488 -193 492
rect -173 488 -169 492
rect -188 454 -184 458
rect -165 454 -161 458
rect -147 487 -143 491
rect -129 488 -125 492
rect -104 488 -100 492
rect -79 487 -75 491
rect 1662 490 1666 494
rect 1718 491 1722 495
rect 82 482 86 486
rect 1990 511 1994 515
rect 1975 477 1979 481
rect 1998 477 2002 481
rect 2016 510 2020 514
rect 2034 511 2038 515
rect 2059 511 2063 515
rect 2084 510 2088 514
rect 2043 477 2047 481
rect 2068 477 2072 481
rect -120 454 -116 458
rect -95 454 -91 458
rect 883 459 887 463
rect 883 451 887 455
rect 77 394 81 398
rect 77 372 81 376
rect 59 362 63 366
rect 884 367 888 371
rect 1680 372 1684 376
rect 115 363 119 367
rect -203 348 -199 352
rect -179 348 -175 352
rect -194 314 -190 318
rect -171 314 -167 318
rect -153 347 -149 351
rect -135 348 -131 352
rect -110 348 -106 352
rect -85 347 -81 351
rect 884 359 888 363
rect 1966 364 1970 368
rect 884 351 888 355
rect 1201 352 1205 356
rect 1201 344 1205 348
rect 1680 350 1684 354
rect 1201 336 1205 340
rect 1662 340 1666 344
rect 1718 341 1722 345
rect 1990 364 1994 368
rect 1975 330 1979 334
rect 1998 330 2002 334
rect 2016 363 2020 367
rect 2034 364 2038 368
rect 2059 364 2063 368
rect 2084 363 2088 367
rect 2043 330 2047 334
rect 2068 330 2072 334
rect -126 314 -122 318
rect -101 314 -97 318
rect 50 307 54 311
rect 50 299 54 303
rect 884 296 888 300
rect 884 288 888 292
rect -203 265 -199 269
rect -179 265 -175 269
rect -194 231 -190 235
rect -171 231 -167 235
rect -153 264 -149 268
rect -135 265 -131 269
rect -110 265 -106 269
rect -85 264 -81 268
rect 82 266 86 270
rect -126 231 -122 235
rect -101 231 -97 235
rect 1680 234 1684 238
rect 882 213 886 217
rect 882 205 886 209
rect 1198 212 1202 216
rect 1967 217 1971 221
rect 1198 204 1202 208
rect 1680 212 1684 216
rect 1662 202 1666 206
rect 1718 203 1722 207
rect 1991 217 1995 221
rect 1976 183 1980 187
rect 1999 183 2003 187
rect 2017 216 2021 220
rect 2035 217 2039 221
rect 2060 217 2064 221
rect 2085 216 2089 220
rect 2044 183 2048 187
rect 2069 183 2073 187
rect 77 178 81 182
rect 77 156 81 160
rect 59 146 63 150
rect 115 147 119 151
rect -216 135 -212 139
rect -192 135 -188 139
rect -207 101 -203 105
rect -184 101 -180 105
rect -166 134 -162 138
rect -148 135 -144 139
rect -123 135 -119 139
rect -98 134 -94 138
rect -139 101 -135 105
rect -114 101 -110 105
rect 1967 112 1971 116
rect 50 91 54 95
rect 50 83 54 87
rect 1991 112 1995 116
rect 1976 78 1980 82
rect 1999 78 2003 82
rect 2017 111 2021 115
rect 2035 112 2039 116
rect 2060 112 2064 116
rect 2085 111 2089 115
rect 2044 78 2048 82
rect 2069 78 2073 82
rect -216 52 -212 56
rect -192 52 -188 56
rect -207 18 -203 22
rect -184 18 -180 22
rect -166 51 -162 55
rect -148 52 -144 56
rect -123 52 -119 56
rect -98 51 -94 55
rect 82 50 86 54
rect -139 18 -135 22
rect -114 18 -110 22
<< metal1 >>
rect 252 1125 1542 1130
rect 236 1117 1525 1122
rect 222 1105 1510 1110
rect 199 1097 202 1102
rect 207 1097 1494 1102
rect 190 1089 1477 1094
rect -73 1066 122 1071
rect -73 1036 -68 1066
rect 58 1051 61 1060
rect 117 1059 122 1066
rect 67 1053 72 1054
rect 117 1054 152 1059
rect 40 1048 61 1051
rect 70 1050 88 1053
rect 58 1045 61 1048
rect 117 1046 120 1054
rect 147 1051 152 1054
rect 147 1046 1741 1051
rect 78 1038 81 1042
rect 108 1041 115 1045
rect -435 1033 -66 1036
rect 40 1035 108 1038
rect 40 1034 43 1035
rect -199 1026 -196 1033
rect -175 1026 -172 1033
rect -149 1026 -146 1033
rect -131 1026 -128 1033
rect -106 1026 -103 1033
rect -81 1026 -78 1033
rect 31 1031 43 1034
rect -242 995 -198 998
rect -182 998 -179 1006
rect -190 995 -174 998
rect -158 998 -155 1006
rect -119 1006 -110 1009
rect -94 1006 -85 1009
rect -141 998 -137 1006
rect -166 995 -148 998
rect -190 994 -187 995
rect -166 994 -163 995
rect -141 995 -130 998
rect -113 998 -110 1006
rect -113 995 -105 998
rect -88 998 -85 1006
rect -73 998 -69 1006
rect -88 995 -80 998
rect -141 990 -137 995
rect -113 994 -110 995
rect -88 994 -85 995
rect -73 995 -3 998
rect -73 990 -69 995
rect -199 971 -196 974
rect -175 971 -172 974
rect -149 971 -146 980
rect -81 974 -78 980
rect -131 971 -128 974
rect -106 971 -103 974
rect -81 971 -35 974
rect -385 968 -78 971
rect -6 972 -3 995
rect -6 969 21 972
rect -343 961 -189 964
rect -185 961 -166 964
rect -162 961 -121 964
rect -117 961 -96 964
rect -7 957 24 960
rect -435 950 -66 953
rect -199 943 -196 950
rect -175 943 -172 950
rect -149 943 -146 950
rect -131 943 -128 950
rect -106 943 -103 950
rect -81 943 -78 950
rect -243 912 -198 915
rect -182 915 -179 923
rect -190 912 -174 915
rect -158 915 -155 923
rect -119 923 -110 926
rect -94 923 -85 926
rect -141 915 -137 923
rect -166 912 -148 915
rect -190 911 -187 912
rect -166 911 -163 912
rect -141 912 -130 915
rect -113 915 -110 923
rect -113 912 -105 915
rect -88 915 -85 923
rect -73 915 -69 923
rect -7 915 -4 957
rect 0 956 24 957
rect 20 951 24 956
rect 31 951 34 1031
rect 64 1026 68 1031
rect 105 1030 108 1035
rect 1012 1034 1017 1046
rect 105 1027 118 1030
rect 59 1025 68 1026
rect 41 1022 55 1025
rect 41 974 44 1022
rect 52 1000 55 1022
rect 59 1014 62 1025
rect 77 1024 80 1027
rect 105 1025 108 1027
rect 75 1013 82 1016
rect 87 1013 90 1016
rect 115 1015 118 1027
rect 128 1026 250 1029
rect 75 1005 88 1008
rect 78 1001 81 1005
rect 951 1006 1116 1011
rect 52 997 59 1000
rect 56 993 59 997
rect 79 996 81 1001
rect 78 993 81 996
rect 953 998 957 1006
rect 56 990 81 993
rect 83 978 125 981
rect 41 959 44 969
rect 58 963 62 969
rect 58 959 67 963
rect 121 959 125 978
rect 253 980 615 981
rect 253 977 888 980
rect 950 979 952 983
rect 984 979 986 983
rect 611 975 888 977
rect 41 956 50 959
rect 46 955 50 956
rect 20 947 50 951
rect 58 947 62 959
rect 137 956 340 959
rect 87 951 97 955
rect 93 947 97 951
rect 58 938 67 947
rect 93 943 101 947
rect 61 936 67 938
rect 63 934 75 936
rect 64 933 75 934
rect 93 933 97 943
rect 57 926 60 928
rect 83 929 97 933
rect 57 923 66 926
rect -88 912 -80 915
rect -141 907 -137 912
rect -113 911 -110 912
rect -88 911 -85 912
rect -73 912 -4 915
rect 63 919 66 923
rect 63 916 71 919
rect -73 907 -69 912
rect 63 903 66 916
rect 83 918 86 929
rect 121 924 123 929
rect 120 919 123 924
rect 113 916 123 919
rect 81 907 93 910
rect -199 888 -196 891
rect -175 888 -172 891
rect -149 888 -146 897
rect -131 888 -128 891
rect -106 888 -103 891
rect -81 888 -78 897
rect 83 896 86 907
rect 120 906 123 916
rect 120 900 123 901
rect 137 896 140 956
rect 83 893 140 896
rect -388 885 -78 888
rect 611 884 615 975
rect 635 967 888 972
rect 963 971 964 975
rect 656 959 888 964
rect 984 963 986 967
rect 701 954 888 955
rect 674 950 888 954
rect 963 955 964 959
rect 674 946 739 950
rect 984 947 986 951
rect 874 942 888 947
rect 895 939 900 943
rect 895 928 899 939
rect 963 939 964 943
rect 895 924 1035 928
rect 936 898 1097 903
rect 936 888 940 898
rect 933 884 940 888
rect 965 884 1012 888
rect -343 878 -189 881
rect -185 878 -166 881
rect -162 878 -121 881
rect -117 878 -96 881
rect 611 880 884 884
rect 936 880 940 884
rect -343 877 -196 878
rect 58 835 61 844
rect 67 837 72 838
rect 117 842 120 844
rect 117 839 128 842
rect 40 832 61 835
rect 70 834 88 837
rect 58 829 61 832
rect 117 830 120 839
rect 78 822 81 826
rect 108 825 115 829
rect -436 818 -64 821
rect 40 819 108 822
rect 40 818 43 819
rect -197 811 -194 818
rect -173 811 -170 818
rect -147 811 -144 818
rect -129 811 -126 818
rect -104 811 -101 818
rect -79 811 -76 818
rect 31 815 43 818
rect -256 780 -196 783
rect -180 783 -177 791
rect -188 780 -172 783
rect -156 783 -153 791
rect -117 791 -108 794
rect -92 791 -83 794
rect -139 783 -135 791
rect -164 780 -146 783
rect -188 779 -185 780
rect -164 779 -161 780
rect -139 780 -128 783
rect -111 783 -108 791
rect -111 780 -103 783
rect -86 783 -83 791
rect -71 783 -67 791
rect -86 780 -78 783
rect -139 775 -135 780
rect -111 779 -108 780
rect -86 779 -83 780
rect -71 780 -1 783
rect -71 775 -67 780
rect -197 756 -194 759
rect -173 756 -170 759
rect -147 756 -144 765
rect -129 756 -126 759
rect -104 756 -101 759
rect -79 756 -76 765
rect -387 753 -76 756
rect -4 756 -1 780
rect -4 753 21 756
rect -343 746 -187 749
rect -183 746 -164 749
rect -160 746 -119 749
rect -115 746 -94 749
rect -5 741 24 744
rect -436 735 -64 738
rect -197 728 -194 735
rect -173 728 -170 735
rect -147 728 -144 735
rect -129 728 -126 735
rect -104 728 -101 735
rect -79 728 -76 735
rect -255 697 -196 700
rect -180 700 -177 708
rect -188 697 -172 700
rect -156 700 -153 708
rect -117 708 -108 711
rect -92 708 -83 711
rect -139 700 -135 708
rect -164 697 -146 700
rect -188 696 -185 697
rect -164 696 -161 697
rect -139 697 -128 700
rect -111 700 -108 708
rect -111 697 -103 700
rect -86 700 -83 708
rect -71 700 -67 708
rect -5 700 -2 741
rect 2 740 24 741
rect 20 735 24 740
rect 31 735 34 815
rect 64 810 68 815
rect 105 814 108 819
rect 105 811 118 814
rect 59 809 68 810
rect 41 806 55 809
rect 41 758 44 806
rect 52 784 55 806
rect 59 798 62 809
rect 77 808 80 811
rect 105 809 108 811
rect 75 797 82 800
rect 87 797 90 800
rect 115 799 118 811
rect 128 810 233 813
rect 75 789 88 792
rect 78 785 81 789
rect 611 788 615 880
rect 936 876 945 880
rect 881 875 884 876
rect 656 872 884 875
rect 881 867 884 868
rect 674 864 884 867
rect 936 864 940 876
rect 971 872 975 884
rect 965 868 975 872
rect 936 860 945 864
rect 874 857 884 860
rect 881 856 884 857
rect 971 856 975 868
rect 891 852 893 856
rect 965 852 975 856
rect 891 844 894 852
rect 891 841 1036 844
rect 1092 833 1097 898
rect 1111 841 1116 1006
rect 1432 891 1687 898
rect 1111 836 1183 841
rect 1245 840 1247 844
rect 1279 840 1281 844
rect 1092 828 1183 833
rect 1258 832 1259 836
rect 1050 821 1183 825
rect 1279 824 1281 828
rect 929 820 1183 821
rect 929 818 1056 820
rect 1084 811 1183 816
rect 1258 816 1259 820
rect 918 789 924 793
rect 955 789 964 793
rect 1084 791 1089 811
rect 1279 808 1281 812
rect 52 781 59 784
rect 56 777 59 781
rect 79 780 81 785
rect 78 777 81 780
rect 56 774 81 777
rect 611 785 881 788
rect 924 785 928 789
rect 83 762 125 765
rect 41 743 44 753
rect 58 747 62 753
rect 58 743 67 747
rect 121 743 125 762
rect 41 740 50 743
rect 46 739 50 740
rect 20 731 50 735
rect 58 731 62 743
rect 137 740 322 743
rect 87 735 97 739
rect 93 731 97 735
rect 58 722 67 731
rect 93 727 101 731
rect 61 720 67 722
rect 63 718 75 720
rect 64 717 75 718
rect 93 717 97 727
rect 57 710 60 712
rect 83 713 97 717
rect 57 707 66 710
rect -86 697 -78 700
rect -139 692 -135 697
rect -111 696 -108 697
rect -86 696 -83 697
rect -71 697 -2 700
rect 63 703 66 707
rect 63 700 71 703
rect -71 692 -67 697
rect 63 684 66 700
rect 83 702 86 713
rect 121 708 123 713
rect 120 703 123 708
rect 113 700 123 703
rect 81 691 93 694
rect -197 673 -194 676
rect -173 673 -170 676
rect -147 673 -144 682
rect -129 673 -126 676
rect -104 673 -101 676
rect -79 673 -76 682
rect 83 680 86 691
rect 120 690 123 700
rect 120 684 123 685
rect 137 680 140 740
rect 611 715 615 785
rect 924 781 935 785
rect 657 777 881 780
rect 735 769 881 772
rect 926 769 930 781
rect 960 777 964 789
rect 955 773 964 777
rect 960 771 964 773
rect 926 765 935 769
rect 960 767 1013 771
rect 899 755 903 765
rect 899 751 1034 755
rect 891 727 1013 731
rect 891 719 895 727
rect 954 720 1034 724
rect 891 715 900 719
rect 954 715 958 720
rect 611 711 883 715
rect 692 704 700 705
rect 707 704 883 707
rect 692 703 883 704
rect 891 703 895 715
rect 920 707 930 711
rect 926 703 930 707
rect 692 700 711 703
rect 692 697 700 700
rect 891 699 900 703
rect 926 699 934 703
rect 926 695 930 699
rect 1085 695 1089 791
rect 926 691 1089 695
rect 1102 803 1183 808
rect 1432 814 1439 891
rect 1736 840 1741 1046
rect 1841 933 2102 936
rect 1969 926 1972 933
rect 1993 926 1996 933
rect 2019 926 2022 933
rect 2037 926 2040 933
rect 2062 926 2065 933
rect 2087 926 2090 933
rect 1786 895 1970 898
rect 1986 898 1989 906
rect 1978 895 1994 898
rect 2010 898 2013 906
rect 2049 906 2058 909
rect 2074 906 2083 909
rect 2027 898 2031 906
rect 2002 895 2020 898
rect 1786 894 1810 895
rect 1978 894 1981 895
rect 2002 894 2005 895
rect 2027 895 2038 898
rect 2055 898 2058 906
rect 2055 895 2063 898
rect 2080 898 2083 906
rect 2095 898 2099 906
rect 2080 895 2088 898
rect 1786 891 1803 894
rect 2027 890 2031 895
rect 2055 894 2058 895
rect 2080 894 2083 895
rect 2095 895 2172 898
rect 2095 890 2099 895
rect 1969 871 1972 874
rect 1993 871 1996 874
rect 2019 871 2022 880
rect 2037 871 2040 874
rect 2062 871 2065 874
rect 2087 871 2090 880
rect 1886 868 2090 871
rect 1929 861 1979 864
rect 1983 861 2002 864
rect 2006 861 2047 864
rect 2051 861 2072 864
rect 1838 846 2106 849
rect 1669 824 1672 840
rect 1678 833 1683 834
rect 1728 837 1744 840
rect 1681 830 1699 833
rect 1658 821 1677 824
rect 1728 825 1731 837
rect 1736 836 1744 837
rect 1689 818 1692 822
rect 1719 821 1731 825
rect 1546 815 1719 818
rect 1346 810 1439 814
rect 1432 809 1439 810
rect 1675 806 1679 811
rect 1716 810 1719 815
rect 1716 807 1729 810
rect 1670 805 1679 806
rect 1102 687 1107 803
rect 1190 800 1195 804
rect 1190 792 1194 800
rect 1258 800 1259 804
rect 1670 794 1673 805
rect 1688 804 1691 807
rect 1716 805 1719 807
rect 1686 793 1693 796
rect 1698 793 1701 796
rect 1726 795 1729 807
rect 1686 785 1699 788
rect 1689 781 1692 785
rect 83 677 140 680
rect 345 679 1107 687
rect 1435 776 1685 780
rect 1690 776 1692 781
rect -387 670 -76 673
rect -344 663 -187 666
rect -183 663 -164 666
rect -160 663 -119 666
rect -115 663 -94 666
rect 938 633 1156 637
rect 58 619 61 628
rect 117 627 120 628
rect 67 621 72 622
rect 117 624 127 627
rect 40 616 61 619
rect 70 618 88 621
rect 58 613 61 616
rect 117 614 120 624
rect 938 623 942 633
rect 935 619 942 623
rect 967 619 1013 623
rect 708 616 886 619
rect -436 609 -65 612
rect -198 602 -195 609
rect -174 602 -171 609
rect -148 602 -145 609
rect -130 602 -127 609
rect -105 602 -102 609
rect -80 602 -77 609
rect 78 606 81 610
rect 108 609 115 613
rect 237 615 886 616
rect 938 615 942 619
rect 237 610 598 615
rect 603 611 719 615
rect 938 611 947 615
rect 603 610 699 611
rect 708 610 719 611
rect 40 603 108 606
rect 40 602 43 603
rect 31 599 43 602
rect -255 571 -197 574
rect -181 574 -178 582
rect -189 571 -173 574
rect -157 574 -154 582
rect -118 582 -109 585
rect -93 582 -84 585
rect -140 574 -136 582
rect -165 571 -147 574
rect -189 570 -186 571
rect -165 570 -162 571
rect -140 571 -129 574
rect -112 574 -109 582
rect -112 571 -104 574
rect -87 574 -84 582
rect -72 574 -68 582
rect -87 571 -79 574
rect -140 566 -136 571
rect -112 570 -109 571
rect -87 570 -84 571
rect -72 571 -3 574
rect -72 566 -68 571
rect -198 547 -195 550
rect -174 547 -171 550
rect -148 547 -145 556
rect -130 547 -127 550
rect -105 547 -102 550
rect -80 547 -77 556
rect -386 544 -77 547
rect -342 537 -188 540
rect -184 537 -165 540
rect -161 537 -120 540
rect -116 537 -95 540
rect -6 540 -3 571
rect -6 537 21 540
rect -435 526 -65 529
rect -198 519 -195 526
rect -174 519 -171 526
rect -148 519 -145 526
rect -130 519 -127 526
rect -105 519 -102 526
rect -80 519 -77 526
rect -7 525 24 528
rect -255 488 -197 491
rect -181 491 -178 499
rect -189 488 -173 491
rect -157 491 -154 499
rect -118 499 -109 502
rect -93 499 -84 502
rect -140 491 -136 499
rect -165 488 -147 491
rect -189 487 -186 488
rect -165 487 -162 488
rect -140 488 -129 491
rect -112 491 -109 499
rect -112 488 -104 491
rect -87 491 -84 499
rect -72 491 -68 499
rect -7 491 -4 525
rect 2 524 24 525
rect 20 519 24 524
rect 31 519 34 599
rect 64 594 68 599
rect 105 598 108 603
rect 655 599 706 602
rect 105 595 118 598
rect 59 593 68 594
rect 41 590 55 593
rect 41 542 44 590
rect 52 568 55 590
rect 59 582 62 593
rect 77 592 80 595
rect 105 593 108 595
rect 75 581 82 584
rect 87 581 90 584
rect 115 583 118 595
rect 128 594 218 597
rect 703 590 707 591
rect 671 587 707 590
rect 75 573 88 576
rect 78 569 81 573
rect 52 565 59 568
rect 56 561 59 565
rect 79 564 81 569
rect 78 561 81 564
rect 56 558 81 561
rect 83 546 125 549
rect 41 527 44 537
rect 58 531 62 537
rect 58 527 67 531
rect 121 527 125 546
rect 713 533 719 610
rect 743 608 886 611
rect 743 605 746 608
rect 883 607 886 608
rect 727 602 746 605
rect 753 600 886 603
rect 753 594 756 600
rect 883 599 886 600
rect 938 599 942 611
rect 973 607 977 619
rect 967 603 977 607
rect 727 591 756 594
rect 938 595 947 599
rect 869 592 886 595
rect 883 591 886 592
rect 973 591 977 603
rect 893 587 895 591
rect 967 587 977 591
rect 893 576 896 587
rect 893 573 1035 576
rect 991 546 1099 549
rect 920 534 926 538
rect 957 534 966 538
rect 713 530 883 533
rect 926 530 930 534
rect 41 524 50 527
rect 46 523 50 524
rect 20 515 50 519
rect 58 515 62 527
rect 137 524 307 527
rect 655 524 703 527
rect 87 519 97 523
rect 93 515 97 519
rect 58 506 67 515
rect 93 511 101 515
rect 61 504 67 506
rect 63 502 75 504
rect 64 501 75 502
rect 93 501 97 511
rect 57 494 60 496
rect 83 497 97 501
rect 57 491 66 494
rect -87 488 -79 491
rect -140 483 -136 488
rect -112 487 -109 488
rect -87 487 -84 488
rect -72 488 -4 491
rect -72 483 -68 488
rect 63 487 66 491
rect 63 484 71 487
rect -198 464 -195 467
rect -174 464 -171 467
rect -148 464 -145 473
rect -130 464 -127 467
rect -105 464 -102 467
rect -80 464 -77 473
rect 63 468 66 484
rect 83 486 86 497
rect 121 492 123 497
rect 120 487 123 492
rect 113 484 123 487
rect 81 475 93 478
rect -386 461 -77 464
rect 83 464 86 475
rect 120 474 123 484
rect 120 468 123 469
rect 137 464 140 524
rect 83 461 140 464
rect 713 463 719 530
rect 926 526 937 530
rect 727 522 883 525
rect 879 514 883 517
rect 928 514 932 526
rect 962 522 966 534
rect 1096 529 1099 546
rect 1152 538 1156 633
rect 1244 556 1319 560
rect 1244 542 1248 556
rect 1241 538 1248 542
rect 1273 538 1291 542
rect 1152 534 1192 538
rect 1244 534 1248 538
rect 1244 530 1253 534
rect 1189 529 1192 530
rect 1096 526 1192 529
rect 957 518 966 522
rect 1189 521 1192 522
rect 962 514 1011 518
rect 1065 518 1192 521
rect 1244 518 1248 530
rect 1279 526 1283 538
rect 1273 522 1283 526
rect 928 510 937 514
rect 962 512 966 514
rect 901 503 905 510
rect 901 499 1034 503
rect 891 475 1013 479
rect 891 467 895 475
rect 954 471 958 472
rect 954 467 1034 471
rect 891 463 900 467
rect 954 463 958 467
rect 713 459 883 463
rect -346 454 -188 457
rect -184 454 -165 457
rect -161 454 -120 457
rect -116 454 -95 457
rect 737 448 876 452
rect 879 448 883 455
rect 891 451 895 463
rect 920 455 930 459
rect 926 451 930 455
rect 737 444 883 448
rect 891 447 900 451
rect 926 447 934 451
rect 926 437 930 447
rect 1065 437 1068 518
rect 1244 514 1253 518
rect 1189 513 1192 514
rect 1156 510 1192 513
rect 1279 510 1283 522
rect 926 433 1071 437
rect 1156 426 1159 510
rect 1199 506 1201 510
rect 1273 506 1283 510
rect 1199 502 1202 506
rect 1287 487 1291 538
rect 1315 517 1319 556
rect 1435 517 1439 776
rect 1659 767 1669 772
rect 1666 550 1669 767
rect 1741 565 1744 836
rect 1973 839 1976 846
rect 1997 839 2000 846
rect 2023 839 2026 846
rect 2041 839 2044 846
rect 2066 839 2069 846
rect 2091 839 2094 846
rect 1760 811 1780 813
rect 1760 810 1974 811
rect 1777 808 1974 810
rect 1990 811 1993 819
rect 1982 808 1998 811
rect 2014 811 2017 819
rect 2053 819 2062 822
rect 2078 819 2087 822
rect 2031 811 2035 819
rect 2006 808 2024 811
rect 1982 807 1985 808
rect 2006 807 2009 808
rect 2031 808 2042 811
rect 2059 811 2062 819
rect 2059 808 2067 811
rect 2084 811 2087 819
rect 2099 811 2103 819
rect 2084 808 2092 811
rect 2031 803 2035 808
rect 2059 807 2062 808
rect 2084 807 2087 808
rect 2099 808 2172 811
rect 2099 803 2103 808
rect 1973 784 1976 787
rect 1997 784 2000 787
rect 2023 784 2026 793
rect 2041 784 2044 787
rect 2066 784 2069 787
rect 2091 784 2094 793
rect 1886 781 2094 784
rect 1929 774 1983 777
rect 1987 774 2006 777
rect 2010 774 2051 777
rect 2055 774 2076 777
rect 1661 547 1669 550
rect 1733 562 1744 565
rect 1661 524 1664 547
rect 1733 540 1736 562
rect 1837 549 2098 552
rect 1670 533 1675 534
rect 1720 537 1736 540
rect 1965 542 1968 549
rect 1989 542 1992 549
rect 2015 542 2018 549
rect 2033 542 2036 549
rect 2058 542 2061 549
rect 2083 542 2086 549
rect 1673 530 1691 533
rect 1650 521 1669 524
rect 1720 525 1723 537
rect 1315 513 1439 517
rect 1681 518 1684 522
rect 1711 521 1723 525
rect 1529 515 1711 518
rect 1667 506 1671 511
rect 1708 510 1711 515
rect 1708 507 1721 510
rect 1662 505 1671 506
rect 1662 494 1665 505
rect 1680 504 1683 507
rect 1708 505 1711 507
rect 1678 493 1685 496
rect 1690 493 1693 496
rect 1718 495 1721 507
rect 1678 485 1691 488
rect 1681 481 1684 485
rect 1435 476 1677 480
rect 1682 476 1684 481
rect 328 418 684 426
rect 692 418 1163 426
rect 58 403 61 412
rect 67 405 72 406
rect 117 410 120 412
rect 117 407 128 410
rect 40 400 61 403
rect 70 402 88 405
rect 58 397 61 400
rect 117 398 120 407
rect 78 390 81 394
rect 108 393 115 397
rect -434 386 -71 389
rect 40 387 108 390
rect 40 386 43 387
rect -204 379 -201 386
rect -180 379 -177 386
rect -154 379 -151 386
rect -136 379 -133 386
rect -111 379 -108 386
rect -86 379 -83 386
rect 31 383 43 386
rect -253 348 -203 351
rect -187 351 -184 359
rect -195 348 -179 351
rect -163 351 -160 359
rect -124 359 -115 362
rect -99 359 -90 362
rect -146 351 -142 359
rect -171 348 -153 351
rect -195 347 -192 348
rect -171 347 -168 348
rect -146 348 -135 351
rect -118 351 -115 359
rect -118 348 -110 351
rect -93 351 -90 359
rect -78 351 -74 359
rect -93 348 -85 351
rect -146 343 -142 348
rect -118 347 -115 348
rect -93 347 -90 348
rect -78 348 -3 351
rect -78 343 -74 348
rect -204 324 -201 327
rect -180 324 -177 327
rect -154 324 -151 333
rect -136 324 -133 327
rect -111 324 -108 327
rect -86 324 -83 333
rect -386 321 -83 324
rect -6 325 -3 348
rect -6 324 10 325
rect -6 322 21 324
rect 5 321 21 322
rect -343 314 -194 317
rect -190 314 -171 317
rect -167 314 -126 317
rect -122 314 -101 317
rect 5 311 24 312
rect -4 308 24 311
rect -434 303 -71 306
rect -204 296 -201 303
rect -180 296 -177 303
rect -154 296 -151 303
rect -136 296 -133 303
rect -111 296 -108 303
rect -86 296 -83 303
rect -254 265 -203 268
rect -187 268 -184 276
rect -195 265 -179 268
rect -163 268 -160 276
rect -124 276 -115 279
rect -99 276 -90 279
rect -146 268 -142 276
rect -171 265 -153 268
rect -195 264 -192 265
rect -171 264 -168 265
rect -146 265 -135 268
rect -118 268 -115 276
rect -118 265 -110 268
rect -93 268 -90 276
rect -78 268 -74 276
rect -4 268 -1 308
rect 20 303 24 308
rect 31 303 34 383
rect 64 378 68 383
rect 105 382 108 387
rect 990 385 1168 388
rect 105 379 118 382
rect 59 377 68 378
rect 41 374 55 377
rect 41 326 44 374
rect 52 352 55 374
rect 59 366 62 377
rect 77 376 80 379
rect 105 377 108 379
rect 75 365 82 368
rect 87 365 90 368
rect 115 367 118 379
rect 128 378 201 381
rect 921 371 927 375
rect 958 371 967 375
rect 220 365 651 370
rect 656 367 884 370
rect 927 367 931 371
rect 656 365 825 367
rect 75 357 88 360
rect 78 353 81 357
rect 52 349 59 352
rect 56 345 59 349
rect 79 348 81 353
rect 78 345 81 348
rect 56 342 81 345
rect 83 330 125 333
rect 41 311 44 321
rect 58 315 62 321
rect 58 311 67 315
rect 121 311 125 330
rect 41 308 50 311
rect 46 307 50 308
rect 20 299 50 303
rect 58 299 62 311
rect 137 308 292 311
rect 87 303 97 307
rect 93 299 97 303
rect 58 290 67 299
rect 93 295 101 299
rect 61 288 67 290
rect 63 286 75 288
rect 64 285 75 286
rect 93 285 97 295
rect 57 278 60 280
rect 83 281 97 285
rect 57 275 66 278
rect -93 265 -85 268
rect -146 260 -142 265
rect -118 264 -115 265
rect -93 264 -90 265
rect -78 265 -1 268
rect 63 271 66 275
rect 63 268 71 271
rect -78 260 -74 265
rect 63 252 66 268
rect 83 270 86 281
rect 121 276 123 281
rect 120 271 123 276
rect 113 268 123 271
rect 81 259 93 262
rect -204 241 -201 244
rect -180 241 -177 244
rect -154 241 -151 250
rect -136 241 -133 244
rect -111 241 -108 244
rect -86 241 -83 250
rect 83 248 86 259
rect 120 258 123 268
rect 120 252 123 253
rect 137 248 140 308
rect 747 300 751 365
rect 927 363 938 367
rect 757 359 884 362
rect 757 340 760 359
rect 869 351 884 354
rect 929 351 933 363
rect 963 359 967 371
rect 958 355 967 359
rect 963 353 967 355
rect 1164 355 1168 385
rect 1238 356 1244 360
rect 1275 356 1284 360
rect 929 347 938 351
rect 963 349 1012 353
rect 1164 352 1201 355
rect 1244 352 1248 356
rect 1244 348 1255 352
rect 1050 347 1054 348
rect 902 338 906 347
rect 1049 344 1201 347
rect 902 334 1033 338
rect 892 312 1013 316
rect 892 304 896 312
rect 955 305 1034 309
rect 892 300 901 304
rect 955 300 959 305
rect 747 296 884 300
rect 878 288 884 292
rect 892 288 896 300
rect 921 292 931 296
rect 927 288 931 292
rect 892 284 901 288
rect 927 284 935 288
rect 927 281 931 284
rect 1050 281 1054 344
rect 927 277 1054 281
rect 1178 336 1201 339
rect 1246 336 1250 348
rect 1280 344 1284 356
rect 1275 340 1284 344
rect 1435 345 1439 476
rect 1651 467 1661 472
rect 1658 407 1661 467
rect 1658 399 1664 407
rect 1661 374 1664 399
rect 1733 390 1736 537
rect 1782 513 1966 514
rect 1752 511 1966 513
rect 1982 514 1985 522
rect 1974 511 1990 514
rect 2006 514 2009 522
rect 2045 522 2054 525
rect 2070 522 2079 525
rect 2023 514 2027 522
rect 1998 511 2016 514
rect 1752 510 1785 511
rect 1974 510 1977 511
rect 1998 510 2001 511
rect 2023 511 2034 514
rect 2051 514 2054 522
rect 2051 511 2059 514
rect 2076 514 2079 522
rect 2091 514 2095 522
rect 2076 511 2084 514
rect 1759 509 1785 510
rect 2023 506 2027 511
rect 2051 510 2054 511
rect 2076 510 2079 511
rect 2091 511 2163 514
rect 2091 506 2095 511
rect 1965 487 1968 490
rect 1989 487 1992 490
rect 2015 487 2018 496
rect 2033 487 2036 490
rect 2058 487 2061 490
rect 2083 487 2086 496
rect 1886 484 2086 487
rect 1930 477 1975 480
rect 1979 477 1998 480
rect 2002 477 2043 480
rect 2047 477 2068 480
rect 1839 402 2098 405
rect 1965 395 1968 402
rect 1989 395 1992 402
rect 2015 395 2018 402
rect 2033 395 2036 402
rect 2058 395 2061 402
rect 2083 395 2086 402
rect 1670 383 1675 384
rect 1720 387 1736 390
rect 1673 380 1691 383
rect 1650 371 1669 374
rect 1720 375 1723 387
rect 1681 368 1684 372
rect 1711 371 1723 375
rect 1516 365 1711 368
rect 1312 342 1439 345
rect 1667 356 1671 361
rect 1708 360 1711 365
rect 1708 357 1721 360
rect 1662 355 1671 356
rect 1662 344 1665 355
rect 1680 354 1683 357
rect 1708 355 1711 357
rect 1678 343 1685 346
rect 1690 343 1693 346
rect 1718 345 1721 357
rect 1178 269 1181 336
rect 1246 332 1255 336
rect 1219 327 1223 332
rect 1280 317 1284 340
rect 1678 335 1691 338
rect 1681 331 1684 335
rect 1427 326 1677 330
rect 1682 326 1684 331
rect 313 261 729 269
rect 737 261 1185 269
rect 1178 260 1181 261
rect 83 245 140 248
rect -386 238 -83 241
rect -345 231 -194 234
rect -190 231 -171 234
rect -167 231 -126 234
rect -122 231 -101 234
rect 890 230 1013 234
rect 1039 233 1069 237
rect 890 221 894 230
rect 1065 229 1273 233
rect 953 225 957 226
rect 953 221 1035 225
rect 1100 222 1210 226
rect 890 217 899 221
rect 953 217 957 221
rect 207 206 666 214
rect 674 212 724 214
rect 729 213 882 217
rect 729 212 733 213
rect 674 208 733 212
rect 674 206 724 208
rect 862 205 882 209
rect 890 205 894 217
rect 1100 217 1104 222
rect 1206 220 1210 222
rect 1017 213 1104 217
rect 1151 214 1198 218
rect 1206 216 1215 220
rect 1269 216 1273 229
rect 919 209 929 213
rect 925 205 929 209
rect 58 187 61 196
rect 67 189 72 190
rect 117 193 120 196
rect 117 190 128 193
rect 40 184 61 187
rect 70 186 88 189
rect 58 181 61 184
rect 117 182 120 190
rect -435 173 -84 176
rect 78 174 81 178
rect 108 177 115 181
rect 862 174 866 205
rect 890 201 899 205
rect 925 201 933 205
rect 925 194 929 201
rect 1151 194 1155 214
rect 1194 212 1198 214
rect 925 190 1155 194
rect 1178 204 1198 208
rect 1206 204 1210 216
rect 1427 212 1431 326
rect 1651 317 1661 322
rect 1658 266 1661 317
rect 1658 263 1664 266
rect 1661 236 1664 263
rect 1733 252 1736 387
rect 1787 364 1966 367
rect 1982 367 1985 375
rect 1974 364 1990 367
rect 2006 367 2009 375
rect 2045 375 2054 378
rect 2070 375 2079 378
rect 2023 367 2027 375
rect 1998 364 2016 367
rect 1758 363 1790 364
rect 1974 363 1977 364
rect 1998 363 2001 364
rect 2023 364 2034 367
rect 2051 367 2054 375
rect 2051 364 2059 367
rect 2076 367 2079 375
rect 2091 367 2095 375
rect 2076 364 2084 367
rect 1752 361 1790 363
rect 1752 360 1761 361
rect 2023 359 2027 364
rect 2051 363 2054 364
rect 2076 363 2079 364
rect 2091 364 2145 367
rect 2091 359 2095 364
rect 1965 340 1968 343
rect 1989 340 1992 343
rect 2015 340 2018 349
rect 2033 340 2036 343
rect 2058 340 2061 343
rect 2083 340 2086 349
rect 1887 337 2086 340
rect 1930 330 1975 333
rect 1979 330 1998 333
rect 2002 330 2043 333
rect 2047 330 2068 333
rect 1837 255 2099 258
rect 1670 245 1675 246
rect 1720 249 1736 252
rect 1673 242 1691 245
rect 1650 233 1669 236
rect 1720 237 1723 249
rect 1681 230 1684 234
rect 1711 233 1723 237
rect 1497 227 1711 230
rect 1235 208 1245 212
rect 1283 209 1431 212
rect 1667 218 1671 223
rect 1708 222 1711 227
rect 1708 219 1721 222
rect 1662 217 1671 218
rect 1283 208 1430 209
rect 1241 204 1245 208
rect 1178 174 1182 204
rect 1206 200 1215 204
rect 1241 200 1249 204
rect 1241 194 1245 200
rect 1283 194 1287 208
rect 1662 206 1665 217
rect 1680 216 1683 219
rect 1708 217 1711 219
rect 1678 205 1685 208
rect 1690 205 1693 208
rect 1718 207 1721 219
rect 1678 197 1691 200
rect 1241 190 1287 194
rect 1681 193 1684 197
rect 1423 188 1677 192
rect 1682 188 1684 193
rect -217 166 -214 173
rect -193 166 -190 173
rect -167 166 -164 173
rect -149 166 -146 173
rect -124 166 -121 173
rect -99 166 -96 173
rect 40 171 108 174
rect 40 170 43 171
rect 31 167 43 170
rect -255 135 -216 138
rect -200 138 -197 146
rect -208 135 -192 138
rect -176 138 -173 146
rect -137 146 -128 149
rect -112 146 -103 149
rect -159 138 -155 146
rect -184 135 -166 138
rect -208 134 -205 135
rect -184 134 -181 135
rect -159 135 -148 138
rect -131 138 -128 146
rect -131 135 -123 138
rect -106 138 -103 146
rect -91 138 -87 146
rect -106 135 -98 138
rect -159 130 -155 135
rect -131 134 -128 135
rect -106 134 -103 135
rect -91 135 -7 138
rect -91 130 -87 135
rect -217 111 -214 114
rect -193 111 -190 114
rect -167 111 -164 120
rect -149 111 -146 114
rect -124 111 -121 114
rect -99 111 -96 120
rect -388 108 -96 111
rect -10 109 -7 135
rect -10 108 8 109
rect -10 106 21 108
rect 4 105 21 106
rect -345 101 -207 104
rect -203 101 -184 104
rect -180 101 -139 104
rect -135 101 -114 104
rect -8 93 24 96
rect -437 90 -84 93
rect -217 83 -214 90
rect -193 83 -190 90
rect -167 83 -164 90
rect -149 83 -146 90
rect -124 83 -121 90
rect -99 83 -96 90
rect -253 52 -216 55
rect -200 55 -197 63
rect -208 52 -192 55
rect -176 55 -173 63
rect -137 63 -128 66
rect -112 63 -103 66
rect -159 55 -155 63
rect -184 52 -166 55
rect -208 51 -205 52
rect -184 51 -181 52
rect -159 52 -148 55
rect -131 55 -128 63
rect -131 52 -123 55
rect -106 55 -103 63
rect -91 55 -87 63
rect -8 55 -5 93
rect 4 92 24 93
rect 20 87 24 92
rect 31 87 34 167
rect 64 162 68 167
rect 105 166 108 171
rect 105 163 118 166
rect 59 161 68 162
rect 41 158 55 161
rect 41 110 44 158
rect 52 136 55 158
rect 59 150 62 161
rect 77 160 80 163
rect 105 161 108 163
rect 75 149 82 152
rect 87 149 90 152
rect 115 151 118 163
rect 128 162 185 165
rect 298 173 1183 174
rect 298 168 722 173
rect 727 168 1183 173
rect 298 166 1183 168
rect 75 141 88 144
rect 78 137 81 141
rect 52 133 59 136
rect 56 129 59 133
rect 79 132 81 137
rect 78 129 81 132
rect 56 126 81 129
rect 281 132 724 134
rect 862 132 866 166
rect 1423 132 1427 188
rect 1651 179 1661 184
rect 1658 136 1661 179
rect 1733 174 1736 249
rect 1966 248 1969 255
rect 1990 248 1993 255
rect 2016 248 2019 255
rect 2034 248 2037 255
rect 2059 248 2062 255
rect 2084 248 2087 255
rect 1752 222 1767 225
rect 1764 220 1767 222
rect 1764 217 1967 220
rect 1983 220 1986 228
rect 1975 217 1991 220
rect 2007 220 2010 228
rect 2046 228 2055 231
rect 2071 228 2080 231
rect 2024 220 2028 228
rect 1999 217 2017 220
rect 1975 216 1978 217
rect 1999 216 2002 217
rect 2024 217 2035 220
rect 2052 220 2055 228
rect 2052 217 2060 220
rect 2077 220 2080 228
rect 2092 220 2096 228
rect 2077 217 2085 220
rect 2024 212 2028 217
rect 2052 216 2055 217
rect 2077 216 2080 217
rect 2092 217 2146 220
rect 2092 212 2096 217
rect 1966 193 1969 196
rect 1990 193 1993 196
rect 2016 193 2019 202
rect 2034 193 2037 196
rect 2059 193 2062 196
rect 2084 193 2087 202
rect 1885 190 2087 193
rect 1929 183 1976 186
rect 1980 183 1999 186
rect 2003 183 2044 186
rect 2048 183 2069 186
rect 1733 171 1836 174
rect 1733 167 1736 171
rect 1838 150 2099 153
rect 1966 143 1969 150
rect 1990 143 1993 150
rect 2016 143 2019 150
rect 2034 143 2037 150
rect 2059 143 2062 150
rect 2084 143 2087 150
rect 1658 133 1885 136
rect 281 128 1431 132
rect 281 126 724 128
rect 773 127 777 128
rect 1484 120 1617 127
rect 83 114 150 117
rect 121 113 150 114
rect 41 95 44 105
rect 58 99 62 105
rect 58 95 67 99
rect 121 95 125 113
rect 41 92 50 95
rect 46 91 50 92
rect 20 83 50 87
rect 58 83 62 95
rect 137 92 276 95
rect 1658 95 1661 133
rect 1709 123 1762 127
rect 1709 120 1772 123
rect 1769 115 1772 120
rect 1769 112 1967 115
rect 1983 115 1986 123
rect 1975 112 1991 115
rect 2007 115 2010 123
rect 2046 123 2055 126
rect 2071 123 2080 126
rect 2024 115 2028 123
rect 1999 112 2017 115
rect 1975 111 1978 112
rect 1999 111 2002 112
rect 2024 112 2035 115
rect 2052 115 2055 123
rect 2052 112 2060 115
rect 2077 115 2080 123
rect 2092 115 2096 123
rect 2077 112 2085 115
rect 2024 107 2028 112
rect 2052 111 2055 112
rect 2077 111 2080 112
rect 2092 112 2143 115
rect 2092 107 2096 112
rect 1442 92 1661 95
rect 87 87 97 91
rect 93 83 97 87
rect 58 74 67 83
rect 93 79 101 83
rect 61 72 67 74
rect 63 70 75 72
rect 64 69 75 70
rect 93 69 97 79
rect 57 62 60 64
rect 83 65 97 69
rect 57 59 66 62
rect -106 52 -98 55
rect -159 47 -155 52
rect -131 51 -128 52
rect -106 51 -103 52
rect -91 52 -5 55
rect 63 55 66 59
rect 63 52 71 55
rect -91 47 -87 52
rect -217 28 -214 31
rect -193 28 -190 31
rect -167 28 -164 37
rect -149 28 -146 31
rect -124 28 -121 31
rect -99 28 -96 37
rect 63 36 66 52
rect 83 54 86 65
rect 121 60 123 65
rect 120 55 123 60
rect 113 52 123 55
rect 81 43 93 46
rect 83 32 86 43
rect 120 42 123 52
rect 120 36 123 37
rect 137 32 140 92
rect 1033 35 1039 53
rect 158 34 1120 35
rect 1442 34 1445 92
rect 1966 88 1969 91
rect 1990 88 1993 91
rect 2016 88 2019 97
rect 2034 88 2037 91
rect 2059 88 2062 91
rect 2084 88 2087 97
rect 1889 85 2087 88
rect 1929 78 1976 81
rect 1980 78 1999 81
rect 2003 78 2044 81
rect 2048 78 2069 81
rect 83 29 140 32
rect 158 32 1445 34
rect 155 31 1445 32
rect 155 29 1120 31
rect 155 28 162 29
rect -387 25 -96 28
rect -343 18 -207 21
rect -203 18 -184 21
rect -180 18 -139 21
rect -135 18 -114 21
<< m2contact >>
rect 247 1125 252 1130
rect 1542 1125 1547 1130
rect 231 1117 236 1122
rect 1525 1117 1530 1122
rect 217 1105 222 1110
rect 1510 1105 1515 1110
rect 202 1097 207 1102
rect 1494 1097 1499 1102
rect 185 1089 190 1094
rect 1477 1089 1482 1094
rect -440 1032 -435 1037
rect 67 1054 72 1059
rect 35 1046 40 1051
rect 115 1041 120 1046
rect -390 967 -385 972
rect -35 970 -30 975
rect 21 968 26 973
rect -348 960 -343 965
rect -440 949 -435 954
rect 59 1026 64 1031
rect 82 1012 87 1017
rect 123 1025 128 1030
rect 250 1026 255 1031
rect 1012 1029 1017 1034
rect 953 993 958 998
rect 78 977 83 982
rect 41 969 46 974
rect 248 977 253 982
rect 952 979 957 984
rect 986 978 991 983
rect 340 956 345 961
rect 55 928 60 933
rect 75 932 80 937
rect 116 924 121 929
rect 63 898 68 903
rect -393 885 -388 890
rect 119 901 124 906
rect 630 967 635 972
rect 958 970 963 975
rect 651 959 656 964
rect 986 962 991 967
rect 666 946 674 954
rect 958 954 963 959
rect 869 942 874 947
rect 986 946 991 951
rect 958 938 963 943
rect 1035 924 1040 929
rect 1012 884 1017 889
rect -348 876 -343 881
rect 67 838 72 843
rect 35 830 40 835
rect 128 838 133 843
rect 115 825 120 830
rect -441 817 -436 822
rect -392 753 -387 758
rect 21 752 26 757
rect -348 745 -343 750
rect -441 735 -436 740
rect 59 810 64 815
rect 82 796 87 801
rect 123 809 128 814
rect 233 810 238 815
rect 651 872 656 877
rect 669 864 674 869
rect 869 856 874 861
rect 1036 841 1041 846
rect 1687 891 1694 898
rect 1247 840 1252 845
rect 1281 839 1286 844
rect 1253 831 1258 836
rect 924 817 929 822
rect 1281 823 1286 828
rect 1253 815 1258 820
rect 924 789 929 794
rect 78 761 83 766
rect 41 753 46 758
rect 322 740 327 745
rect 55 712 60 717
rect 75 716 80 721
rect 116 708 121 713
rect -392 670 -387 675
rect 119 685 124 690
rect 652 777 657 782
rect 730 769 735 774
rect 1013 767 1018 772
rect 1034 751 1039 756
rect 1013 727 1018 732
rect 1034 720 1039 725
rect 684 697 692 705
rect 1281 807 1286 812
rect 1341 810 1346 815
rect 1836 932 1841 937
rect 1779 891 1786 898
rect 1881 867 1886 872
rect 1924 860 1929 865
rect 1833 845 1838 850
rect 1653 821 1658 826
rect 1678 834 1683 839
rect 1541 814 1546 819
rect 1670 806 1675 811
rect 1253 799 1258 804
rect 1190 787 1195 792
rect 1693 792 1698 797
rect 337 679 345 687
rect -349 662 -344 667
rect 67 622 72 627
rect 35 614 40 619
rect -441 609 -436 614
rect 127 623 132 628
rect 1013 619 1018 624
rect 115 609 120 614
rect 231 610 237 616
rect 598 610 603 615
rect -391 544 -386 549
rect -347 536 -342 541
rect 21 536 26 541
rect -440 526 -435 531
rect 59 594 64 599
rect 650 599 655 604
rect 701 602 706 607
rect 82 580 87 585
rect 123 593 128 598
rect 218 594 223 599
rect 666 587 671 592
rect 78 545 83 550
rect 41 537 46 542
rect 722 601 727 606
rect 722 591 727 596
rect 864 592 869 597
rect 1035 573 1040 578
rect 986 545 991 550
rect 926 534 931 539
rect 307 524 312 529
rect 650 524 655 529
rect 55 496 60 501
rect 75 500 80 505
rect -391 460 -386 465
rect 116 492 121 497
rect 119 469 124 474
rect 703 523 708 528
rect 722 521 727 526
rect 874 514 879 519
rect 1034 499 1039 504
rect 1013 475 1018 480
rect 1034 467 1039 472
rect -351 453 -346 458
rect 729 444 737 452
rect 1199 497 1204 502
rect 1654 767 1659 772
rect 1755 809 1760 814
rect 1881 780 1886 785
rect 1924 773 1929 778
rect 1645 521 1650 526
rect 1832 549 1837 554
rect 1670 534 1675 539
rect 1524 515 1529 520
rect 1662 506 1667 511
rect 1685 492 1690 497
rect 1287 482 1292 487
rect 320 418 328 426
rect 684 418 692 426
rect 67 406 72 411
rect 35 398 40 403
rect 128 406 133 411
rect -439 386 -434 391
rect 115 393 120 398
rect -391 320 -386 325
rect 21 320 26 325
rect -348 313 -343 318
rect -439 303 -434 308
rect 59 378 64 383
rect 985 384 990 389
rect 82 364 87 369
rect 123 377 128 382
rect 201 378 206 383
rect 927 371 932 376
rect 215 365 220 370
rect 651 365 656 370
rect 78 329 83 334
rect 41 321 46 326
rect 292 308 297 313
rect 55 280 60 285
rect 75 284 80 289
rect 116 276 121 281
rect -391 238 -386 243
rect 119 253 124 258
rect 864 351 869 356
rect 1244 356 1249 361
rect 1012 349 1017 354
rect 756 335 761 340
rect 1013 312 1018 317
rect 1034 305 1039 310
rect 873 288 878 293
rect 1307 341 1312 346
rect 1646 467 1651 472
rect 1645 371 1650 376
rect 1747 509 1752 514
rect 1881 484 1886 489
rect 1925 476 1930 481
rect 1834 401 1839 406
rect 1670 384 1675 389
rect 1511 365 1516 370
rect 1662 356 1667 361
rect 1685 342 1690 347
rect 1219 322 1224 327
rect 1280 312 1285 317
rect 305 261 313 269
rect 729 261 737 269
rect -350 230 -345 235
rect 1013 230 1018 235
rect 1034 233 1039 238
rect 1035 221 1040 226
rect 199 206 207 214
rect 666 206 674 214
rect 1012 213 1017 218
rect 67 190 72 195
rect 35 182 40 187
rect 128 189 133 194
rect -440 173 -435 178
rect 115 177 120 182
rect 1646 317 1651 322
rect 1645 233 1650 238
rect 1747 359 1752 364
rect 1882 337 1887 342
rect 1925 329 1930 334
rect 1832 254 1837 259
rect 1670 246 1675 251
rect 1492 227 1497 232
rect 1662 218 1667 223
rect 1685 204 1690 209
rect -393 108 -388 113
rect -350 100 -345 105
rect 21 104 26 109
rect -442 90 -437 95
rect 59 162 64 167
rect 82 148 87 153
rect 123 161 128 166
rect 185 162 190 167
rect 290 166 298 174
rect 722 168 727 173
rect 273 126 281 134
rect 773 132 778 137
rect 1646 179 1651 184
rect 1747 221 1752 226
rect 1880 189 1885 194
rect 1924 182 1929 187
rect 1836 171 1841 176
rect 1833 150 1838 155
rect 1885 133 1890 138
rect 1477 120 1484 127
rect 1617 120 1624 127
rect 78 113 83 118
rect 150 113 155 118
rect 41 105 46 110
rect 1702 120 1709 127
rect 55 64 60 69
rect 75 68 80 73
rect -392 25 -387 30
rect 116 60 121 65
rect 119 37 124 42
rect 1033 53 1039 59
rect 1884 85 1889 90
rect 1924 77 1929 82
rect 150 28 155 33
rect -348 17 -343 22
<< pdm12contact >>
rect 703 591 708 596
rect 1011 514 1016 519
rect 1033 334 1038 339
rect 276 92 281 97
<< metal2 >>
rect -444 1037 -430 1112
rect -444 1032 -440 1037
rect -435 1032 -430 1037
rect -444 954 -430 1032
rect -444 949 -440 954
rect -435 949 -430 954
rect -444 822 -430 949
rect -444 817 -441 822
rect -436 817 -430 822
rect -444 740 -430 817
rect -444 735 -441 740
rect -436 735 -430 740
rect -444 614 -430 735
rect -444 609 -441 614
rect -436 609 -430 614
rect -444 531 -430 609
rect -444 526 -440 531
rect -435 526 -430 531
rect -444 391 -430 526
rect -444 386 -439 391
rect -434 386 -430 391
rect -444 308 -430 386
rect -444 303 -439 308
rect -434 303 -430 308
rect -444 178 -430 303
rect -444 173 -440 178
rect -435 173 -430 178
rect -444 95 -430 173
rect -444 90 -442 95
rect -437 90 -430 95
rect -444 0 -430 90
rect -396 972 -382 1110
rect -396 967 -390 972
rect -385 967 -382 972
rect -396 890 -382 967
rect -396 885 -393 890
rect -388 885 -382 890
rect -396 758 -382 885
rect -396 753 -392 758
rect -387 753 -382 758
rect -396 675 -382 753
rect -396 670 -392 675
rect -387 670 -382 675
rect -396 549 -382 670
rect -396 544 -391 549
rect -386 544 -382 549
rect -396 465 -382 544
rect -396 460 -391 465
rect -386 460 -382 465
rect -396 325 -382 460
rect -396 320 -391 325
rect -386 320 -382 325
rect -396 243 -382 320
rect -396 238 -391 243
rect -386 238 -382 243
rect -396 113 -382 238
rect -396 108 -393 113
rect -388 108 -382 113
rect -396 30 -382 108
rect -396 25 -392 30
rect -387 25 -382 30
rect -396 0 -382 25
rect -354 965 -340 1110
rect 184 1094 191 1134
rect 184 1089 185 1094
rect 190 1089 191 1094
rect 46 1055 67 1058
rect -35 1047 25 1050
rect -35 975 -32 1047
rect 30 1047 35 1050
rect 46 1031 49 1055
rect 116 1040 120 1041
rect 46 1028 59 1031
rect 83 994 86 1012
rect 123 994 126 1025
rect 83 991 126 994
rect 73 979 78 982
rect 26 970 41 973
rect -354 960 -348 965
rect -343 960 -340 965
rect -354 881 -340 960
rect 75 928 78 932
rect 75 925 116 928
rect 126 927 130 933
rect 126 924 131 927
rect -354 876 -348 881
rect -343 876 -340 881
rect -354 750 -340 876
rect -354 745 -348 750
rect -343 745 -340 750
rect -354 667 -340 745
rect -354 662 -349 667
rect -344 662 -340 667
rect -354 541 -340 662
rect -354 536 -347 541
rect -342 536 -340 541
rect -354 458 -340 536
rect 14 899 63 902
rect 14 717 17 899
rect 128 905 131 924
rect 124 902 131 905
rect 128 843 131 902
rect 46 839 67 842
rect 30 831 35 834
rect 46 815 49 839
rect 116 824 120 825
rect 46 812 59 815
rect 83 778 86 796
rect 123 778 126 809
rect 83 775 126 778
rect 73 763 78 766
rect 26 754 41 757
rect 184 750 191 1089
rect 183 743 191 750
rect 14 714 55 717
rect 14 500 17 714
rect 75 712 78 716
rect 75 709 116 712
rect 126 711 130 717
rect 126 708 131 711
rect 128 689 131 708
rect 124 686 131 689
rect 128 628 131 686
rect 46 623 67 626
rect 30 615 35 618
rect 46 599 49 623
rect 116 608 120 609
rect 46 596 59 599
rect 83 562 86 580
rect 123 562 126 593
rect 83 559 126 562
rect 73 547 78 550
rect 26 538 41 541
rect 10 497 55 500
rect -354 453 -351 458
rect -346 453 -340 458
rect -354 318 -340 453
rect -354 313 -348 318
rect -343 313 -340 318
rect -354 235 -340 313
rect -354 230 -350 235
rect -345 230 -340 235
rect -354 105 -340 230
rect -354 100 -350 105
rect -345 100 -340 105
rect -354 22 -340 100
rect 13 284 16 497
rect 75 496 78 500
rect 75 493 116 496
rect 126 495 130 501
rect 126 492 131 495
rect 184 494 191 743
rect 128 473 131 492
rect 183 487 191 494
rect 124 470 131 473
rect 128 411 131 470
rect 46 407 67 410
rect 30 399 35 402
rect 46 383 49 407
rect 116 392 120 393
rect 46 380 59 383
rect 83 346 86 364
rect 123 346 126 377
rect 83 343 126 346
rect 73 331 78 334
rect 26 322 41 325
rect 13 281 55 284
rect 13 69 16 281
rect 75 280 78 284
rect 75 277 116 280
rect 126 279 130 285
rect 126 276 131 279
rect 128 257 131 276
rect 124 254 131 257
rect 46 191 67 194
rect 30 183 35 186
rect 46 167 49 191
rect 128 194 131 254
rect 184 195 191 487
rect 183 188 191 195
rect 116 176 120 177
rect 46 164 59 167
rect 184 167 191 188
rect 184 162 185 167
rect 190 162 191 167
rect 83 130 86 148
rect 123 130 126 161
rect 83 127 126 130
rect 73 115 78 118
rect 26 106 41 109
rect 13 66 55 69
rect 75 64 78 68
rect 75 61 116 64
rect 126 63 130 69
rect 126 60 131 63
rect 128 41 131 60
rect 124 38 131 41
rect 150 33 154 113
rect -354 17 -348 22
rect -343 17 -340 22
rect -354 -110 -340 17
rect 184 2 191 162
rect 199 1102 206 1134
rect 216 1110 223 1135
rect 216 1105 217 1110
rect 222 1105 223 1110
rect 199 1097 202 1102
rect 199 750 206 1097
rect 216 750 223 1105
rect 231 1122 238 1136
rect 236 1117 238 1122
rect 231 815 238 1117
rect 231 810 233 815
rect 231 750 238 810
rect 247 1130 254 1135
rect 252 1125 254 1130
rect 247 1031 254 1125
rect 247 1026 250 1031
rect 247 982 254 1026
rect 247 977 248 982
rect 253 977 254 982
rect 247 750 254 977
rect 274 750 281 1136
rect 290 750 297 1136
rect 199 743 207 750
rect 215 743 223 750
rect 230 743 238 750
rect 246 743 254 750
rect 273 743 281 750
rect 289 743 297 750
rect 199 494 206 743
rect 216 599 223 743
rect 216 594 218 599
rect 216 494 223 594
rect 231 616 238 743
rect 237 610 238 616
rect 231 494 238 610
rect 247 494 254 743
rect 274 494 281 743
rect 290 494 297 743
rect 199 487 207 494
rect 215 487 223 494
rect 230 487 238 494
rect 246 487 254 494
rect 273 487 281 494
rect 289 487 297 494
rect 199 383 206 487
rect 199 378 201 383
rect 199 214 206 378
rect 216 370 223 487
rect 220 365 223 370
rect 199 195 206 206
rect 216 195 223 365
rect 231 195 238 487
rect 247 195 254 487
rect 274 195 281 487
rect 290 313 297 487
rect 290 308 292 313
rect 290 195 297 308
rect 199 188 207 195
rect 215 188 223 195
rect 230 188 238 195
rect 246 188 254 195
rect 273 188 281 195
rect 289 188 297 195
rect 199 2 206 188
rect 216 2 223 188
rect 231 3 238 188
rect 247 0 254 188
rect 274 134 281 188
rect 274 97 281 126
rect 274 92 276 97
rect 274 0 281 92
rect 290 174 297 188
rect 305 750 312 1136
rect 320 750 327 1135
rect 337 961 344 1136
rect 1477 1094 1484 1161
rect 1482 1089 1484 1094
rect 953 984 957 993
rect 1012 983 1017 1029
rect 953 975 957 979
rect 991 979 1017 983
rect 598 967 630 972
rect 953 971 958 975
rect 337 956 340 961
rect 337 750 344 956
rect 305 743 313 750
rect 320 745 328 750
rect 305 529 312 743
rect 305 524 307 529
rect 305 494 312 524
rect 320 740 322 745
rect 327 743 328 745
rect 336 743 344 750
rect 320 494 327 740
rect 337 687 344 743
rect 337 494 344 679
rect 598 615 603 967
rect 651 877 656 959
rect 958 959 962 970
rect 986 967 990 978
rect 651 782 656 872
rect 666 869 674 946
rect 855 942 869 947
rect 958 943 962 954
rect 986 951 990 962
rect 666 864 669 869
rect 651 777 652 782
rect 651 604 656 777
rect 655 599 656 604
rect 651 529 656 599
rect 655 524 656 529
rect 305 487 313 494
rect 320 487 328 494
rect 336 487 344 494
rect 305 269 312 487
rect 320 426 327 487
rect 305 195 312 261
rect 320 195 327 418
rect 337 195 344 487
rect 651 370 656 524
rect 666 592 674 864
rect 1012 889 1017 979
rect 766 860 869 861
rect 765 858 869 860
rect 671 587 674 592
rect 666 346 674 587
rect 684 426 692 697
rect 706 603 722 606
rect 708 592 722 595
rect 708 523 722 526
rect 731 452 734 769
rect 765 518 769 858
rect 924 797 927 817
rect 923 794 927 797
rect 1012 783 1017 884
rect 1033 929 1039 995
rect 1033 924 1035 929
rect 1033 846 1039 924
rect 1248 859 1345 863
rect 1033 841 1036 846
rect 1248 845 1252 859
rect 1033 791 1039 841
rect 1248 836 1252 840
rect 1286 840 1295 844
rect 1248 832 1253 836
rect 1253 820 1257 831
rect 1281 828 1285 839
rect 1253 804 1257 815
rect 1281 812 1285 823
rect 1033 787 1190 791
rect 1012 780 1027 783
rect 1012 779 1023 780
rect 1012 772 1017 779
rect 1012 767 1013 772
rect 1012 732 1017 767
rect 1033 756 1039 787
rect 1291 779 1295 840
rect 1341 815 1345 859
rect 1137 775 1295 779
rect 1033 751 1034 756
rect 1012 727 1013 732
rect 1012 624 1017 727
rect 1033 725 1039 751
rect 1033 720 1034 725
rect 1012 619 1013 624
rect 860 593 864 596
rect 926 545 986 548
rect 926 542 929 545
rect 925 539 929 542
rect 1012 519 1017 619
rect 765 515 874 518
rect 711 348 712 350
rect 729 352 737 444
rect 717 349 754 352
rect 711 346 717 348
rect 665 343 717 346
rect 666 340 717 343
rect 666 214 674 340
rect 729 269 737 349
rect 755 340 758 348
rect 755 336 756 340
rect 765 292 769 515
rect 1016 514 1017 519
rect 1012 490 1017 514
rect 1033 578 1039 720
rect 1033 573 1035 578
rect 1033 504 1039 573
rect 1033 499 1034 504
rect 1039 499 1199 501
rect 1033 498 1199 499
rect 1012 487 1026 490
rect 1012 486 1022 487
rect 1012 480 1017 486
rect 1012 475 1013 480
rect 927 384 985 387
rect 927 379 930 384
rect 926 376 930 379
rect 860 352 864 355
rect 1012 354 1017 475
rect 1012 317 1017 349
rect 1033 472 1039 498
rect 1093 482 1287 486
rect 1033 467 1034 472
rect 1033 339 1039 467
rect 1243 373 1310 376
rect 1243 364 1246 373
rect 1243 361 1247 364
rect 1307 346 1310 373
rect 1038 334 1039 339
rect 1033 326 1039 334
rect 1033 322 1219 326
rect 1012 312 1013 317
rect 1018 312 1023 316
rect 750 288 873 292
rect 305 188 313 195
rect 320 188 328 195
rect 336 188 344 195
rect 290 0 297 166
rect 305 1 312 188
rect 320 2 327 188
rect 337 2 344 188
rect 750 172 754 288
rect 1012 235 1017 312
rect 1033 310 1039 322
rect 1117 312 1280 316
rect 1033 305 1034 310
rect 1033 238 1039 305
rect 1012 230 1013 235
rect 1033 233 1034 238
rect 1012 218 1017 230
rect 1012 185 1017 213
rect 1033 226 1039 233
rect 1033 221 1035 226
rect 727 168 754 172
rect 773 137 777 144
rect 1033 59 1039 221
rect 1477 127 1484 1089
rect 1477 15 1484 120
rect 1492 1102 1499 1163
rect 1492 1097 1494 1102
rect 1492 232 1499 1097
rect 1497 227 1499 232
rect 1492 15 1499 227
rect 1509 1110 1516 1164
rect 1509 1105 1510 1110
rect 1515 1105 1516 1110
rect 1509 370 1516 1105
rect 1509 365 1511 370
rect 1509 15 1516 365
rect 1524 1122 1531 1164
rect 1524 1117 1525 1122
rect 1530 1117 1531 1122
rect 1524 520 1531 1117
rect 1529 515 1531 520
rect 1524 15 1531 515
rect 1540 1130 1547 1163
rect 1540 1125 1542 1130
rect 1540 819 1547 1125
rect 1829 937 1843 1121
rect 1829 932 1836 937
rect 1841 932 1843 937
rect 1694 891 1779 898
rect 1829 850 1843 932
rect 1829 845 1833 850
rect 1838 845 1843 850
rect 1665 835 1678 838
rect 1540 814 1541 819
rect 1546 814 1547 819
rect 1540 15 1547 814
rect 1654 772 1657 821
rect 1665 811 1668 835
rect 1665 808 1670 811
rect 1735 809 1755 812
rect 1694 776 1697 792
rect 1735 776 1738 809
rect 1694 773 1738 776
rect 1829 554 1843 845
rect 1829 549 1832 554
rect 1837 549 1843 554
rect 1657 535 1670 538
rect 1646 472 1649 521
rect 1657 511 1660 535
rect 1657 508 1662 511
rect 1727 509 1747 512
rect 1686 476 1689 492
rect 1727 476 1730 509
rect 1686 473 1730 476
rect 1829 406 1843 549
rect 1829 401 1834 406
rect 1839 401 1843 406
rect 1657 385 1670 388
rect 1646 322 1649 371
rect 1657 361 1660 385
rect 1657 358 1662 361
rect 1727 359 1747 362
rect 1686 326 1689 342
rect 1727 326 1730 359
rect 1686 323 1730 326
rect 1829 259 1843 401
rect 1829 254 1832 259
rect 1837 254 1843 259
rect 1657 247 1670 250
rect 1646 184 1649 233
rect 1657 223 1660 247
rect 1657 220 1662 223
rect 1727 221 1747 224
rect 1686 188 1689 204
rect 1727 188 1730 221
rect 1686 185 1730 188
rect 1829 176 1843 254
rect 1829 171 1836 176
rect 1841 171 1843 176
rect 1829 155 1843 171
rect 1829 150 1833 155
rect 1838 150 1843 155
rect 1624 120 1702 127
rect 1829 77 1843 150
rect 1877 872 1891 1119
rect 1877 867 1881 872
rect 1886 867 1891 872
rect 1877 785 1891 867
rect 1877 780 1881 785
rect 1886 780 1891 785
rect 1877 489 1891 780
rect 1877 484 1881 489
rect 1886 484 1891 489
rect 1877 342 1891 484
rect 1877 337 1882 342
rect 1887 337 1891 342
rect 1877 194 1891 337
rect 1877 189 1880 194
rect 1885 189 1891 194
rect 1877 138 1891 189
rect 1877 133 1885 138
rect 1890 133 1891 138
rect 1877 90 1891 133
rect 1877 85 1884 90
rect 1889 85 1891 90
rect 1877 77 1891 85
rect 1919 865 1933 1119
rect 1919 860 1924 865
rect 1929 860 1933 865
rect 1919 778 1933 860
rect 1919 773 1924 778
rect 1929 773 1933 778
rect 1919 481 1933 773
rect 1919 476 1925 481
rect 1930 476 1933 481
rect 1919 334 1933 476
rect 1919 329 1925 334
rect 1930 329 1933 334
rect 1919 187 1933 329
rect 1919 182 1924 187
rect 1929 182 1933 187
rect 1919 82 1933 182
rect 1919 77 1924 82
rect 1929 77 1933 82
rect 1919 -110 1933 77
rect -354 -124 1936 -110
rect 1919 -125 1933 -124
<< m3contact >>
rect 25 1046 30 1051
rect 116 1035 121 1040
rect 68 978 73 983
rect 60 928 65 933
rect 126 933 131 938
rect 25 830 30 835
rect 116 819 121 824
rect 68 762 73 767
rect 60 712 65 717
rect 126 717 131 722
rect 25 614 30 619
rect 116 603 121 608
rect 68 546 73 551
rect 60 496 65 501
rect 126 501 131 506
rect 25 398 30 403
rect 116 387 121 392
rect 68 330 73 335
rect 60 280 65 285
rect 126 285 131 290
rect 25 182 30 187
rect 116 171 121 176
rect 68 114 73 119
rect 60 64 65 69
rect 126 69 131 74
rect 850 942 855 947
rect 1023 775 1028 780
rect 1132 775 1137 780
rect 855 592 860 597
rect 712 348 717 353
rect 754 348 759 353
rect 1022 482 1027 487
rect 855 351 860 356
rect 1088 482 1093 487
rect 1023 312 1028 317
rect 1112 312 1117 317
rect 773 144 778 149
<< m123contact >>
rect 76 1027 81 1032
rect 74 996 79 1001
rect 76 811 81 816
rect 74 780 79 785
rect 76 595 81 600
rect 74 564 79 569
rect 76 379 81 384
rect 74 348 79 353
rect 76 163 81 168
rect 74 132 79 137
rect 1687 807 1692 812
rect 1685 776 1690 781
rect 1679 507 1684 512
rect 1677 476 1682 481
rect 1679 357 1684 362
rect 1677 326 1682 331
rect 1679 219 1684 224
rect 1677 188 1682 193
<< metal3 >>
rect 24 1051 31 1052
rect 24 1046 25 1051
rect 30 1046 31 1051
rect 24 1045 31 1046
rect 27 1038 30 1045
rect 35 1040 64 1043
rect 35 1038 39 1040
rect 27 1035 39 1038
rect 61 984 64 1040
rect 115 1040 122 1041
rect 115 1035 116 1040
rect 121 1035 122 1040
rect 115 1034 122 1035
rect 77 1001 80 1027
rect 79 998 80 1001
rect 61 983 74 984
rect 61 978 68 983
rect 73 978 74 983
rect 61 977 74 978
rect 61 934 64 977
rect 116 938 120 1034
rect 849 947 856 948
rect 773 942 850 947
rect 855 942 856 947
rect 125 938 132 939
rect 116 934 126 938
rect 59 933 65 934
rect 125 933 126 934
rect 131 933 132 938
rect 59 928 60 933
rect 65 928 66 933
rect 125 932 132 933
rect 59 927 66 928
rect 24 835 31 836
rect 24 830 25 835
rect 30 830 31 835
rect 24 829 31 830
rect 27 822 30 829
rect 35 824 64 827
rect 35 822 39 824
rect 27 819 39 822
rect 61 768 64 824
rect 115 824 122 825
rect 115 819 116 824
rect 121 819 122 824
rect 115 818 122 819
rect 77 785 80 811
rect 79 782 80 785
rect 61 767 74 768
rect 61 762 68 767
rect 73 762 74 767
rect 61 761 74 762
rect 61 718 64 761
rect 116 722 120 818
rect 125 722 132 723
rect 116 718 126 722
rect 59 717 65 718
rect 125 717 126 718
rect 131 717 132 722
rect 59 712 60 717
rect 65 712 66 717
rect 125 716 132 717
rect 59 711 66 712
rect 24 619 31 620
rect 24 614 25 619
rect 30 614 31 619
rect 24 613 31 614
rect 27 606 30 613
rect 35 608 64 611
rect 35 606 39 608
rect 27 603 39 606
rect 61 552 64 608
rect 115 608 122 609
rect 115 603 116 608
rect 121 603 122 608
rect 115 602 122 603
rect 77 569 80 595
rect 79 566 80 569
rect 61 551 74 552
rect 61 546 68 551
rect 73 546 74 551
rect 61 545 74 546
rect 61 502 64 545
rect 116 506 120 602
rect 774 596 778 942
rect 849 941 856 942
rect 1688 781 1691 807
rect 1022 780 1029 781
rect 1022 775 1023 780
rect 1028 779 1029 780
rect 1131 780 1138 781
rect 1131 779 1132 780
rect 1028 775 1132 779
rect 1137 775 1138 780
rect 1690 778 1691 781
rect 1022 774 1029 775
rect 1131 774 1138 775
rect 854 597 861 598
rect 854 596 855 597
rect 774 593 855 596
rect 125 506 132 507
rect 116 502 126 506
rect 59 501 65 502
rect 125 501 126 502
rect 131 501 132 506
rect 59 496 60 501
rect 65 496 66 501
rect 125 500 132 501
rect 59 495 66 496
rect 24 403 31 404
rect 24 398 25 403
rect 30 398 31 403
rect 24 397 31 398
rect 27 390 30 397
rect 35 392 64 395
rect 35 390 39 392
rect 27 387 39 390
rect 61 336 64 392
rect 115 392 122 393
rect 115 387 116 392
rect 121 387 122 392
rect 115 386 122 387
rect 77 353 80 379
rect 79 350 80 353
rect 61 335 74 336
rect 61 330 68 335
rect 73 330 74 335
rect 61 329 74 330
rect 61 286 64 329
rect 116 290 120 386
rect 774 355 778 593
rect 854 592 855 593
rect 860 592 861 597
rect 854 591 861 592
rect 1021 487 1028 488
rect 1021 482 1022 487
rect 1027 486 1028 487
rect 1087 487 1094 488
rect 1087 486 1088 487
rect 1027 482 1088 486
rect 1093 482 1094 487
rect 1021 481 1028 482
rect 1087 481 1094 482
rect 1680 481 1683 507
rect 1682 478 1683 481
rect 854 356 861 357
rect 854 355 855 356
rect 711 353 718 354
rect 711 348 712 353
rect 717 352 718 353
rect 753 353 760 354
rect 753 352 754 353
rect 717 349 754 352
rect 717 348 718 349
rect 711 347 718 348
rect 753 348 754 349
rect 759 348 760 353
rect 753 347 760 348
rect 774 352 855 355
rect 125 290 132 291
rect 116 286 126 290
rect 59 285 65 286
rect 125 285 126 286
rect 131 285 132 290
rect 59 280 60 285
rect 65 280 66 285
rect 125 284 132 285
rect 59 279 66 280
rect 24 187 31 188
rect 24 182 25 187
rect 30 182 31 187
rect 24 181 31 182
rect 27 174 30 181
rect 35 176 64 179
rect 35 174 39 176
rect 27 171 39 174
rect 61 120 64 176
rect 115 176 122 177
rect 115 171 116 176
rect 121 171 122 176
rect 115 170 122 171
rect 77 137 80 163
rect 79 134 80 137
rect 61 119 74 120
rect 61 114 68 119
rect 73 114 74 119
rect 61 113 74 114
rect 61 70 64 113
rect 116 74 120 170
rect 774 150 778 352
rect 854 351 855 352
rect 860 351 861 356
rect 854 350 861 351
rect 1680 331 1683 357
rect 1682 328 1683 331
rect 1022 317 1029 318
rect 1022 312 1023 317
rect 1028 316 1029 317
rect 1111 317 1118 318
rect 1111 316 1112 317
rect 1028 312 1112 316
rect 1117 312 1118 317
rect 1022 311 1029 312
rect 1111 311 1118 312
rect 1680 193 1683 219
rect 1682 190 1683 193
rect 772 149 779 150
rect 772 144 773 149
rect 778 144 779 149
rect 772 143 779 144
rect 125 74 132 75
rect 116 70 126 74
rect 59 69 65 70
rect 125 69 126 70
rect 131 69 132 74
rect 59 64 60 69
rect 65 64 66 69
rect 125 68 132 69
rect 59 63 66 64
<< labels >>
rlabel metal1 64 918 64 918 3 gnd
rlabel metal1 64 702 64 702 3 gnd
rlabel metal1 64 486 64 486 3 gnd
rlabel metal1 64 270 64 270 3 gnd
rlabel metal1 64 54 64 54 3 gnd
rlabel metal1 122 919 122 919 7 vdd
rlabel metal1 122 703 122 703 7 vdd
rlabel metal1 122 487 122 487 7 vdd
rlabel metal1 122 271 122 271 7 vdd
rlabel metal1 122 55 122 55 7 vdd
rlabel metal1 46 947 54 951 3 input_1
port 1 s
rlabel metal1 46 731 54 735 3 input_2
port 1 s
rlabel metal1 46 515 54 519 3 input_3
port 1 s
rlabel metal1 46 299 54 303 3 input_4
port 1 s
rlabel metal1 46 83 54 87 3 input_5
port 1 s
rlabel metal1 46 955 54 959 3 input_2
port 2 s
rlabel metal1 46 739 54 743 3 input_3
port 2 s
rlabel metal1 46 523 54 527 3 input_4
port 2 s
rlabel metal1 46 307 54 311 3 input_5
port 2 s
rlabel metal1 46 91 54 95 3 input_6
port 2 s
rlabel metal1 121 959 125 968 7 ground
port 5 n
rlabel metal1 121 743 125 752 7 ground
port 5 n
rlabel metal1 121 527 125 536 7 ground
port 5 n
rlabel metal1 121 311 125 320 7 ground
port 5 n
rlabel metal1 121 95 125 104 7 ground
port 5 n
rlabel metal1 58 960 62 969 5 power_supply
port 3 w
rlabel metal1 58 744 62 753 5 power_supply
port 3 w
rlabel metal1 58 528 62 537 5 power_supply
port 3 w
rlabel metal1 58 312 62 321 5 power_supply
port 3 w
rlabel metal1 58 96 62 105 5 power_supply
port 3 w
rlabel metal1 93 939 97 943 1 output
port 4 e
rlabel metal1 93 723 97 727 1 output
port 4 e
rlabel metal1 93 507 97 511 1 output
port 4 e
rlabel metal1 93 291 97 295 1 output
port 4 e
rlabel metal1 93 75 97 79 1 output
port 4 e
rlabel metal1 118 1054 118 1054 7 vdd
rlabel metal1 118 838 118 838 7 vdd
rlabel metal1 118 622 118 622 7 vdd
rlabel metal1 118 406 118 406 7 vdd
rlabel metal1 118 190 118 190 7 vdd
rlabel metal1 78 1035 80 1038 1 in1
rlabel metal1 78 819 80 822 1 in2
rlabel metal1 78 603 80 606 1 in3
rlabel metal1 78 387 80 390 1 in4
rlabel metal1 78 171 80 174 1 in5
rlabel m2contact 60 1029 60 1029 3 in1_inv
rlabel m2contact 60 813 60 813 3 in2_inv
rlabel m2contact 60 597 60 597 3 in3_inv
rlabel m2contact 60 381 60 381 3 in4_inv
rlabel m2contact 60 165 60 165 3 in5_inv
rlabel metal3 80 1003 80 1003 3 in2
rlabel metal3 80 787 80 787 3 in3
rlabel metal3 80 571 80 571 3 in4
rlabel metal3 80 355 80 355 3 in5
rlabel metal3 80 139 80 139 3 in6
rlabel space 476 113 495 139 1 G0
rlabel space 480 156 499 182 1 G1
rlabel space 480 200 499 226 1 P1
rlabel space 479 250 498 276 1 G2
rlabel space 473 356 492 382 1 P2
rlabel space 479 406 498 432 1 G3
rlabel space 471 598 490 624 1 P3
rlabel space 474 667 493 693 1 G4
rlabel space 460 967 479 993 1 P4
rlabel space 1411 115 1440 141 1 C1
rlabel space 1410 197 1439 223 1 C2
rlabel space 1418 329 1447 355 1 C3
rlabel space 1419 502 1448 528 1 C4
rlabel space 1418 798 1447 824 1 C5
rlabel space 450 21 479 47 1 ground
rlabel space 471 1036 500 1062 5 power
rlabel metal1 1684 495 1684 495 3 out
rlabel metal3 1683 483 1683 483 3 in2
rlabel m2contact 1663 509 1663 509 3 in1_inv
rlabel metal1 1681 515 1683 518 1 in1
rlabel metal1 1662 525 1662 525 3 gnd
rlabel metal1 1721 534 1721 534 7 vdd
rlabel metal1 1684 345 1684 345 3 out
rlabel metal3 1683 333 1683 333 3 in2
rlabel m2contact 1663 359 1663 359 3 in1_inv
rlabel metal1 1681 365 1683 368 1 in1
rlabel metal1 1662 375 1662 375 3 gnd
rlabel metal1 1721 384 1721 384 7 vdd
rlabel metal1 1684 207 1684 207 3 out
rlabel metal3 1683 195 1683 195 3 in2
rlabel m2contact 1663 221 1663 221 3 in1_inv
rlabel metal1 1681 227 1683 230 1 in1
rlabel metal1 1662 237 1662 237 3 gnd
rlabel metal1 1721 246 1721 246 7 vdd
rlabel metal1 1692 795 1692 795 3 out
rlabel metal3 1691 783 1691 783 3 in2
rlabel m2contact 1671 809 1671 809 3 in1_inv
rlabel metal1 1689 815 1691 818 1 in1
rlabel metal1 1670 825 1670 825 3 gnd
rlabel metal1 1729 834 1729 834 7 vdd
rlabel metal1 -222 54 -222 54 1 d
rlabel metal1 -216 91 -216 91 5 vdd
rlabel metal1 -221 19 -221 19 1 clk
rlabel metal1 -198 26 -198 26 1 gnd
rlabel metal1 -86 53 -86 53 7 q
rlabel metal1 -222 137 -222 137 1 d
rlabel metal1 -216 174 -216 174 5 vdd
rlabel metal1 -221 102 -221 102 1 clk
rlabel metal1 -198 109 -198 109 1 gnd
rlabel metal1 -86 136 -86 136 7 q
rlabel metal1 -209 267 -209 267 1 d
rlabel metal1 -203 304 -203 304 5 vdd
rlabel metal1 -208 232 -208 232 1 clk
rlabel metal1 -185 239 -185 239 1 gnd
rlabel metal1 -73 266 -73 266 7 q
rlabel metal1 -209 350 -209 350 1 d
rlabel metal1 -203 387 -203 387 5 vdd
rlabel metal1 -208 315 -208 315 1 clk
rlabel metal1 -185 322 -185 322 1 gnd
rlabel metal1 -73 349 -73 349 7 q
rlabel metal1 -203 490 -203 490 1 d
rlabel metal1 -197 527 -197 527 5 vdd
rlabel metal1 -202 455 -202 455 1 clk
rlabel metal1 -179 462 -179 462 1 gnd
rlabel metal1 -67 489 -67 489 7 q
rlabel metal1 -203 573 -203 573 1 d
rlabel metal1 -197 610 -197 610 5 vdd
rlabel metal1 -202 538 -202 538 1 clk
rlabel metal1 -179 545 -179 545 1 gnd
rlabel metal1 -67 572 -67 572 7 q
rlabel metal1 -202 699 -202 699 1 d
rlabel metal1 -196 736 -196 736 5 vdd
rlabel metal1 -201 664 -201 664 1 clk
rlabel metal1 -178 671 -178 671 1 gnd
rlabel metal1 -66 698 -66 698 7 q
rlabel metal1 -202 782 -202 782 1 d
rlabel metal1 -196 819 -196 819 5 vdd
rlabel metal1 -201 747 -201 747 1 clk
rlabel metal1 -178 754 -178 754 1 gnd
rlabel metal1 -66 781 -66 781 7 q
rlabel metal1 -68 996 -68 996 7 q
rlabel metal1 -180 969 -180 969 1 gnd
rlabel metal1 -203 962 -203 962 1 clk
rlabel metal1 -198 1034 -198 1034 5 vdd
rlabel metal1 -204 997 -204 997 1 d
rlabel metal1 -68 913 -68 913 7 q
rlabel metal1 -180 886 -180 886 1 gnd
rlabel metal1 -203 879 -203 879 1 clk
rlabel metal1 -198 951 -198 951 5 vdd
rlabel metal1 -204 914 -204 914 1 d
rlabel metal1 2104 809 2104 809 7 q
rlabel metal1 1992 782 1992 782 1 gnd
rlabel metal1 1969 775 1969 775 1 clk
rlabel metal1 1974 847 1974 847 5 vdd
rlabel metal1 1968 810 1968 810 1 d
rlabel metal1 2096 512 2096 512 7 q
rlabel metal1 1984 485 1984 485 1 gnd
rlabel metal1 1961 478 1961 478 1 clk
rlabel metal1 1966 550 1966 550 5 vdd
rlabel metal1 1960 513 1960 513 1 d
rlabel metal1 2096 365 2096 365 7 q
rlabel metal1 1984 338 1984 338 1 gnd
rlabel metal1 1961 331 1961 331 1 clk
rlabel metal1 1966 403 1966 403 5 vdd
rlabel metal1 1960 366 1960 366 1 d
rlabel metal1 2097 218 2097 218 7 q
rlabel metal1 1985 191 1985 191 1 gnd
rlabel metal1 1962 184 1962 184 1 clk
rlabel metal1 1967 256 1967 256 5 vdd
rlabel metal1 1961 219 1961 219 1 d
rlabel metal1 2097 113 2097 113 7 q
rlabel metal1 1985 86 1985 86 1 gnd
rlabel metal1 1962 79 1962 79 1 clk
rlabel metal1 1967 151 1967 151 5 vdd
rlabel metal1 1961 114 1961 114 1 d
rlabel metal1 1964 897 1964 897 1 d
rlabel metal1 1970 934 1970 934 5 vdd
rlabel metal1 1965 862 1965 862 1 clk
rlabel metal1 1988 869 1988 869 1 gnd
rlabel metal1 2100 896 2100 896 7 q
rlabel metal1 -253 52 -249 55 1 A1
rlabel metal1 -255 135 -251 138 1 B1
rlabel metal1 -254 265 -250 268 1 A2
rlabel metal1 -253 348 -249 351 1 B2
rlabel metal1 -255 488 -251 491 1 A3
rlabel metal1 -255 571 -251 574 1 B3
rlabel metal1 -255 697 -251 700 1 A4
rlabel metal1 -256 780 -252 783 1 B4
rlabel metal1 -243 912 -239 915 1 A5
rlabel metal1 -242 995 -238 998 1 B5
rlabel metal1 2139 112 2143 115 1 S1
rlabel metal1 2142 217 2146 220 1 S2
rlabel metal1 2141 364 2145 367 1 S3
rlabel metal1 2159 511 2163 514 1 S4
rlabel metal1 2168 808 2172 811 7 S5
rlabel metal1 2168 895 2172 898 7 Cout
<< end >>
