magic
tech scmos
timestamp 1764431408
<< nwell >>
rect -6 26 17 27
rect -6 -5 26 26
<< ntransistor >>
rect 5 -33 7 -13
rect 13 -33 15 -13
<< ptransistor >>
rect 5 1 7 21
rect 13 1 15 21
<< ndiffusion >>
rect 4 -33 5 -13
rect 7 -33 8 -13
rect 12 -33 13 -13
rect 15 -33 16 -13
<< pdiffusion >>
rect 4 1 5 21
rect 7 1 8 21
rect 12 1 13 21
rect 15 1 16 21
<< ndcontact >>
rect 0 -33 4 -13
rect 8 -33 12 -13
rect 16 -33 20 -13
<< pdcontact >>
rect 0 1 4 21
rect 8 1 12 21
rect 16 1 20 21
<< polysilicon >>
rect 5 21 7 34
rect 13 21 15 34
rect 5 -13 7 1
rect 13 -13 15 1
rect 5 -38 7 -33
rect 13 -38 15 -33
<< polycontact >>
rect 4 34 8 38
rect 12 34 16 38
<< metal1 >>
rect 4 38 8 42
rect 12 38 16 42
rect 0 26 26 30
rect 0 21 4 26
rect 16 21 20 26
rect 8 -5 12 1
rect -4 -9 12 -5
rect 0 -13 4 -9
rect 16 -37 25 -33
<< labels >>
rlabel metal1 4 34 8 42 5 input_1
port 1 s
rlabel metal1 12 34 16 42 5 input_2
port 2 s
rlabel metal1 16 -37 25 -33 1 ground
port 5 n
rlabel metal1 17 26 26 30 7 power_supply
port 3 w
rlabel metal1 -4 -9 0 -5 3 output
port 4 e
<< end >>
