.include TSMC_180nm.txt

.param SUPPLY=1.8
.global gnd vdd

VDD vdd gnd SUPPLY
vinA A gnd PULSE(0 SUPPLY   10ns 1ps 1ps   10ns  20ns)
vinB B gnd PULSE(0 SUPPLY    5ns 1ps 1ps    5ns  10ns)
vinC C gnd PULSE(0 SUPPLY  2.5ns 1ps 1ps  2.5ns   5ns)
vinD D gnd PULSE(0 SUPPLY 1.25ns 1ps 1ps 1.25ns 2.5ns)

.option scale=90n

M1000 gnd D a_1_n57# Gnd CMOSN w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=46u
M1001 vdd B output w_n28_n11# CMOSP w=20 l=2
+  ad=60p pd=26u as=60p ps=26u
M1002 vdd D output w_n28_n11# CMOSP w=20 l=2
+  ad=100p pd=50u as=60p ps=26u
M1003 output C vdd w_n28_n11# CMOSP w=20 l=2
+  ad=60p pd=26u as=60p ps=26u
M1004 output A vdd w_n28_n11# CMOSP w=20 l=2
+  ad=60p pd=26u as=100p ps=50u
M1005 a_n7_n57# B a_n15_n57# Gnd CMOSN w=40 l=2
+  ad=0.12n pd=46u as=0.12n ps=46u
M1006 a_1_n57# C a_n7_n57# Gnd CMOSN w=40 l=2
+  ad=0.12n pd=46u as=0.12n ps=46u
M1007 a_n15_n57# A output Gnd CMOSN w=40 l=2
+  ad=0.12n pd=46u as=0.2n ps=90u
C0 vdd A 0.00145f
C1 A w_n28_n11# 0.01842f
C2 B vdd 0.00145f
C3 output C 0.00849f
C4 B w_n28_n11# 0.01803f
C5 vdd output 0.94582f
C6 B A 0.17037f
C7 output w_n28_n11# 0.02246f
C8 D C 0.17037f
C9 a_n15_n57# output 0.46742f
C10 a_n15_n57# a_n7_n57# 0.41238f
C11 output A 0.0097f
C12 vdd D 0.00145f
C13 B output 0.00865f
C14 D w_n28_n11# 0.01842f
C15 gnd a_1_n57# 0.41238f
C16 vdd C 0.00145f
C17 a_n7_n57# output 0.05504f
C18 w_n28_n11# C 0.01803f
C19 D gnd 0
C20 output a_1_n57# 0.05501f
C21 a_n7_n57# a_1_n57# 0.41238f
C22 vdd w_n28_n11# 0.02419f
C23 D output 0.00234f
C24 B C 0.17037f
C25 gnd 0 0.06411f 
C26 a_1_n57# 0 0.00535f 
C27 a_n7_n57# 0 0.00535f 
C28 a_n15_n57# 0 0.00535f 
C29 output 0 0.15501f 
C30 vdd 0 0.19544f 
C31 D 0 0.13691f 
C32 C 0 0.08746f 
C33 B 0 0.08746f 
C34 A 0 0.14017f 
C35 w_n28_n11# 0 1.54276f 


.tran 1n 20n 

.control
  run
  set curplottitle="2024102023_4_NAND"
  * Plot output, and inputs shifted for visibility
  plot  v(A) v(B)+3 v(C)+6 v(D)+9 v(output)+12
.endc

.end