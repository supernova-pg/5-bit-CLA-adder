magic
tech scmos
timestamp 1731385397
<< nwell >>
rect 110 2 252 34
<< ntransistor >>
rect 121 -24 123 -4
rect 145 -24 147 -4
rect 171 -18 173 -8
rect 189 -24 191 -4
rect 198 -24 200 -4
rect 214 -24 216 -4
rect 223 -24 225 -4
rect 239 -18 241 -8
<< ptransistor >>
rect 121 8 123 28
rect 129 8 131 28
rect 145 8 147 28
rect 153 8 155 28
rect 171 8 173 28
rect 189 8 191 28
rect 214 8 216 28
rect 239 8 241 28
<< ndiffusion >>
rect 116 -20 121 -4
rect 120 -24 121 -20
rect 123 -8 124 -4
rect 123 -24 128 -8
rect 140 -20 145 -4
rect 144 -24 145 -20
rect 147 -8 148 -4
rect 147 -24 152 -8
rect 166 -14 171 -8
rect 170 -18 171 -14
rect 173 -12 174 -8
rect 173 -18 178 -12
rect 184 -20 189 -4
rect 188 -24 189 -20
rect 191 -24 198 -4
rect 200 -8 201 -4
rect 200 -24 205 -8
rect 209 -20 214 -4
rect 213 -24 214 -20
rect 216 -24 223 -4
rect 225 -8 226 -4
rect 225 -24 230 -8
rect 234 -14 239 -8
rect 238 -18 239 -14
rect 241 -12 242 -8
rect 241 -18 246 -12
<< pdiffusion >>
rect 120 24 121 28
rect 116 8 121 24
rect 123 8 129 28
rect 131 12 136 28
rect 131 8 132 12
rect 144 24 145 28
rect 140 8 145 24
rect 147 8 153 28
rect 155 12 160 28
rect 155 8 156 12
rect 170 24 171 28
rect 166 8 171 24
rect 173 12 178 28
rect 173 8 174 12
rect 188 24 189 28
rect 184 8 189 24
rect 191 12 196 28
rect 191 8 192 12
rect 213 24 214 28
rect 209 8 214 24
rect 216 12 221 28
rect 216 8 217 12
rect 238 24 239 28
rect 234 8 239 24
rect 241 12 246 28
rect 241 8 242 12
<< ndcontact >>
rect 116 -24 120 -20
rect 124 -8 128 -4
rect 140 -24 144 -20
rect 148 -8 152 -4
rect 166 -18 170 -14
rect 174 -12 178 -8
rect 184 -24 188 -20
rect 201 -8 205 -4
rect 209 -24 213 -20
rect 226 -8 230 -4
rect 234 -18 238 -14
rect 242 -12 246 -8
<< pdcontact >>
rect 116 24 120 28
rect 132 8 136 12
rect 140 24 144 28
rect 156 8 160 12
rect 166 24 170 28
rect 174 8 178 12
rect 184 24 188 28
rect 192 8 196 12
rect 209 24 213 28
rect 217 8 221 12
rect 234 24 238 28
rect 242 8 246 12
<< polysilicon >>
rect 121 28 123 32
rect 129 28 131 32
rect 145 28 147 32
rect 153 28 155 32
rect 171 28 173 32
rect 189 28 191 31
rect 214 28 216 31
rect 239 28 241 32
rect 121 -4 123 8
rect 121 -27 123 -24
rect 129 -33 131 8
rect 145 -4 147 8
rect 145 -27 147 -24
rect 130 -36 131 -33
rect 153 -36 155 8
rect 171 -8 173 8
rect 189 -4 191 8
rect 198 -4 200 0
rect 214 -4 216 8
rect 223 -4 225 0
rect 171 -22 173 -18
rect 239 -8 241 8
rect 239 -22 241 -18
rect 189 -29 191 -24
rect 198 -38 200 -24
rect 214 -29 216 -24
rect 223 -38 225 -24
<< polycontact >>
rect 117 -3 121 1
rect 141 -3 145 1
rect 126 -37 130 -33
rect 149 -37 153 -33
rect 167 -4 171 0
rect 185 -3 189 1
rect 210 -3 214 1
rect 235 -4 239 0
rect 194 -37 198 -33
rect 219 -37 223 -33
<< metal1 >>
rect 116 35 249 38
rect 116 28 119 35
rect 140 28 143 35
rect 166 28 169 35
rect 184 28 187 35
rect 209 28 212 35
rect 234 28 237 35
rect 110 -3 117 0
rect 133 0 136 8
rect 125 -3 141 0
rect 157 0 160 8
rect 196 8 205 11
rect 221 8 230 11
rect 174 0 178 8
rect 149 -3 167 0
rect 125 -4 128 -3
rect 149 -4 152 -3
rect 174 -3 185 0
rect 202 0 205 8
rect 202 -3 210 0
rect 227 0 230 8
rect 242 0 246 8
rect 227 -3 235 0
rect 174 -8 178 -3
rect 202 -4 205 -3
rect 227 -4 230 -3
rect 242 -3 249 0
rect 242 -8 246 -3
rect 116 -27 119 -24
rect 140 -27 143 -24
rect 166 -27 169 -18
rect 184 -27 187 -24
rect 209 -27 212 -24
rect 234 -27 237 -18
rect 116 -30 237 -27
rect 110 -37 126 -34
rect 130 -37 149 -34
rect 153 -37 194 -34
rect 198 -37 219 -34
<< labels >>
rlabel metal1 111 -1 111 -1 1 d
rlabel metal1 117 36 117 36 5 vdd
rlabel metal1 112 -36 112 -36 1 clk
rlabel metal1 135 -29 135 -29 1 gnd
rlabel metal1 247 -2 247 -2 7 q
<< end >>
