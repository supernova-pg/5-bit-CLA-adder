magic
tech scmos
timestamp 1764693657
<< nwell >>
rect 75 732 107 788
rect 56 645 88 693
rect 46 558 78 598
rect 370 593 402 649
rect 11 492 43 524
rect 58 380 90 428
rect 48 303 80 343
rect 364 299 396 347
rect 11 240 43 272
rect 49 140 81 180
rect 366 125 398 165
rect 12 77 44 109
rect 10 -6 42 26
rect 326 -7 358 25
<< ntransistor >>
rect 17 775 67 777
rect 17 767 67 769
rect 17 759 67 761
rect 17 751 67 753
rect 17 743 67 745
rect 10 680 50 682
rect 10 672 50 674
rect 10 664 50 666
rect 10 656 50 658
rect 312 636 362 638
rect 312 628 362 630
rect 312 620 362 622
rect 312 612 362 614
rect 312 604 362 606
rect 5 585 35 587
rect 5 577 35 579
rect 5 569 35 571
rect 51 511 71 513
rect 51 503 71 505
rect 12 415 52 417
rect 12 407 52 409
rect 12 399 52 401
rect 12 391 52 393
rect 318 334 358 336
rect 7 330 37 332
rect 318 326 358 328
rect 7 322 37 324
rect 7 314 37 316
rect 318 318 358 320
rect 318 310 358 312
rect 51 259 71 261
rect 51 251 71 253
rect 8 167 38 169
rect 8 159 38 161
rect 8 151 38 153
rect 325 152 355 154
rect 325 144 355 146
rect 325 136 355 138
rect 52 96 72 98
rect 52 88 72 90
rect 50 13 70 15
rect 366 12 386 14
rect 50 5 70 7
rect 366 4 386 6
<< ptransistor >>
rect 81 775 101 777
rect 81 767 101 769
rect 81 759 101 761
rect 81 751 101 753
rect 81 743 101 745
rect 62 680 82 682
rect 62 672 82 674
rect 62 664 82 666
rect 62 656 82 658
rect 376 636 396 638
rect 376 628 396 630
rect 376 620 396 622
rect 376 612 396 614
rect 376 604 396 606
rect 52 585 72 587
rect 52 577 72 579
rect 52 569 72 571
rect 17 511 37 513
rect 17 503 37 505
rect 64 415 84 417
rect 64 407 84 409
rect 64 399 84 401
rect 64 391 84 393
rect 370 334 390 336
rect 54 330 74 332
rect 370 326 390 328
rect 54 322 74 324
rect 54 314 74 316
rect 370 318 390 320
rect 370 310 390 312
rect 17 259 37 261
rect 17 251 37 253
rect 55 167 75 169
rect 55 159 75 161
rect 55 151 75 153
rect 372 152 392 154
rect 372 144 392 146
rect 372 136 392 138
rect 18 96 38 98
rect 18 88 38 90
rect 16 13 36 15
rect 332 12 352 14
rect 16 5 36 7
rect 332 4 352 6
<< ndiffusion >>
rect 17 777 67 778
rect 17 774 67 775
rect 17 769 67 770
rect 17 766 67 767
rect 17 761 67 762
rect 17 758 67 759
rect 17 753 67 754
rect 17 750 67 751
rect 17 745 67 746
rect 17 742 67 743
rect 10 682 50 683
rect 10 679 50 680
rect 10 674 50 675
rect 10 671 50 672
rect 10 666 50 667
rect 10 663 50 664
rect 10 658 50 659
rect 10 655 50 656
rect 312 638 362 639
rect 312 635 362 636
rect 312 630 362 631
rect 312 627 362 628
rect 312 622 362 623
rect 312 619 362 620
rect 312 614 362 615
rect 312 611 362 612
rect 312 606 362 607
rect 312 603 362 604
rect 5 587 35 588
rect 5 584 35 585
rect 5 579 35 580
rect 5 576 35 577
rect 5 571 35 572
rect 5 568 35 569
rect 51 513 71 514
rect 51 510 71 511
rect 51 505 71 506
rect 51 502 71 503
rect 12 417 52 418
rect 12 414 52 415
rect 12 409 52 410
rect 12 406 52 407
rect 12 401 52 402
rect 12 398 52 399
rect 12 393 52 394
rect 12 390 52 391
rect 7 332 37 333
rect 318 336 358 337
rect 318 333 358 334
rect 7 329 37 330
rect 7 324 37 325
rect 318 328 358 329
rect 318 325 358 326
rect 7 321 37 322
rect 7 316 37 317
rect 7 313 37 314
rect 318 320 358 321
rect 318 317 358 318
rect 318 312 358 313
rect 318 309 358 310
rect 51 261 71 262
rect 51 258 71 259
rect 51 253 71 254
rect 51 250 71 251
rect 8 169 38 170
rect 8 166 38 167
rect 8 161 38 162
rect 8 158 38 159
rect 8 153 38 154
rect 325 154 355 155
rect 325 151 355 152
rect 8 150 38 151
rect 325 146 355 147
rect 325 143 355 144
rect 325 138 355 139
rect 325 135 355 136
rect 52 98 72 99
rect 52 95 72 96
rect 52 90 72 91
rect 52 87 72 88
rect 50 15 70 16
rect 50 12 70 13
rect 366 14 386 15
rect 50 7 70 8
rect 50 4 70 5
rect 366 11 386 12
rect 366 6 386 7
rect 366 3 386 4
<< pdiffusion >>
rect 81 777 101 778
rect 81 774 101 775
rect 81 769 101 770
rect 81 766 101 767
rect 81 761 101 762
rect 81 758 101 759
rect 81 753 101 754
rect 81 750 101 751
rect 81 745 101 746
rect 81 742 101 743
rect 62 682 82 683
rect 62 679 82 680
rect 62 674 82 675
rect 62 671 82 672
rect 62 666 82 667
rect 62 663 82 664
rect 62 658 82 659
rect 62 655 82 656
rect 376 638 396 639
rect 376 635 396 636
rect 376 630 396 631
rect 376 627 396 628
rect 376 622 396 623
rect 376 619 396 620
rect 376 614 396 615
rect 376 611 396 612
rect 376 606 396 607
rect 376 603 396 604
rect 52 587 72 588
rect 52 584 72 585
rect 52 579 72 580
rect 52 576 72 577
rect 52 571 72 572
rect 52 568 72 569
rect 17 513 37 514
rect 17 510 37 511
rect 17 505 37 506
rect 17 502 37 503
rect 64 417 84 418
rect 64 414 84 415
rect 64 409 84 410
rect 64 406 84 407
rect 64 401 84 402
rect 64 398 84 399
rect 64 393 84 394
rect 64 390 84 391
rect 370 336 390 337
rect 54 332 74 333
rect 54 329 74 330
rect 370 333 390 334
rect 370 328 390 329
rect 54 324 74 325
rect 54 321 74 322
rect 54 316 74 317
rect 54 313 74 314
rect 370 325 390 326
rect 370 320 390 321
rect 370 317 390 318
rect 370 312 390 313
rect 370 309 390 310
rect 17 261 37 262
rect 17 258 37 259
rect 17 253 37 254
rect 17 250 37 251
rect 55 169 75 170
rect 55 166 75 167
rect 55 161 75 162
rect 55 158 75 159
rect 55 153 75 154
rect 372 154 392 155
rect 55 150 75 151
rect 372 151 392 152
rect 372 146 392 147
rect 372 143 392 144
rect 372 138 392 139
rect 372 135 392 136
rect 18 98 38 99
rect 18 95 38 96
rect 18 90 38 91
rect 18 87 38 88
rect 16 15 36 16
rect 16 12 36 13
rect 16 7 36 8
rect 332 14 352 15
rect 332 11 352 12
rect 16 4 36 5
rect 332 6 352 7
rect 332 3 352 4
<< ndcontact >>
rect 17 778 67 782
rect 17 770 67 774
rect 17 762 67 766
rect 17 754 67 758
rect 17 746 67 750
rect 17 738 67 742
rect 10 683 50 687
rect 10 675 50 679
rect 10 667 50 671
rect 10 659 50 663
rect 10 651 50 655
rect 312 639 362 643
rect 312 631 362 635
rect 312 623 362 627
rect 312 615 362 619
rect 312 607 362 611
rect 312 599 362 603
rect 5 588 35 592
rect 5 580 35 584
rect 5 572 35 576
rect 5 564 35 568
rect 51 514 71 518
rect 51 506 71 510
rect 51 498 71 502
rect 12 418 52 422
rect 12 410 52 414
rect 12 402 52 406
rect 12 394 52 398
rect 12 386 52 390
rect 318 337 358 341
rect 7 333 37 337
rect 7 325 37 329
rect 318 329 358 333
rect 7 317 37 321
rect 318 321 358 325
rect 7 309 37 313
rect 318 313 358 317
rect 318 305 358 309
rect 51 262 71 266
rect 51 254 71 258
rect 51 246 71 250
rect 8 170 38 174
rect 8 162 38 166
rect 8 154 38 158
rect 325 155 355 159
rect 8 146 38 150
rect 325 147 355 151
rect 325 139 355 143
rect 325 131 355 135
rect 52 99 72 103
rect 52 91 72 95
rect 52 83 72 87
rect 50 16 70 20
rect 50 8 70 12
rect 366 15 386 19
rect 50 0 70 4
rect 366 7 386 11
rect 366 -1 386 3
<< pdcontact >>
rect 81 778 101 782
rect 81 770 101 774
rect 81 762 101 766
rect 81 754 101 758
rect 81 746 101 750
rect 81 738 101 742
rect 62 683 82 687
rect 62 675 82 679
rect 62 667 82 671
rect 62 659 82 663
rect 62 651 82 655
rect 376 639 396 643
rect 376 631 396 635
rect 376 623 396 627
rect 376 615 396 619
rect 376 607 396 611
rect 376 599 396 603
rect 52 588 72 592
rect 52 580 72 584
rect 52 572 72 576
rect 52 564 72 568
rect 17 514 37 518
rect 17 506 37 510
rect 17 498 37 502
rect 64 418 84 422
rect 64 410 84 414
rect 64 402 84 406
rect 64 394 84 398
rect 64 386 84 390
rect 54 333 74 337
rect 370 337 390 341
rect 54 325 74 329
rect 370 329 390 333
rect 54 317 74 321
rect 370 321 390 325
rect 54 309 74 313
rect 370 313 390 317
rect 370 305 390 309
rect 17 262 37 266
rect 17 254 37 258
rect 17 246 37 250
rect 55 170 75 174
rect 55 162 75 166
rect 55 154 75 158
rect 372 155 392 159
rect 55 146 75 150
rect 372 147 392 151
rect 372 139 392 143
rect 372 131 392 135
rect 18 99 38 103
rect 18 91 38 95
rect 18 83 38 87
rect 16 16 36 20
rect 332 15 352 19
rect 16 8 36 12
rect 332 7 352 11
rect 16 0 36 4
rect 332 -1 352 3
<< polysilicon >>
rect 9 775 17 777
rect 67 775 81 777
rect 101 775 104 777
rect 9 767 17 769
rect 67 767 81 769
rect 101 767 104 769
rect 9 759 17 761
rect 67 759 81 761
rect 101 759 104 761
rect 9 751 17 753
rect 67 751 81 753
rect 101 751 104 753
rect 9 743 17 745
rect 67 743 81 745
rect 101 743 104 745
rect 5 680 10 682
rect 50 680 62 682
rect 82 680 85 682
rect 5 672 10 674
rect 50 672 62 674
rect 82 672 85 674
rect 5 664 10 666
rect 50 664 62 666
rect 82 664 85 666
rect 5 656 10 658
rect 50 656 62 658
rect 82 656 85 658
rect 304 636 312 638
rect 362 636 376 638
rect 396 636 399 638
rect 304 628 312 630
rect 362 628 376 630
rect 396 628 399 630
rect 304 620 312 622
rect 362 620 376 622
rect 396 620 399 622
rect 304 612 312 614
rect 362 612 376 614
rect 396 612 399 614
rect 304 604 312 606
rect 362 604 376 606
rect 396 604 399 606
rect 2 585 5 587
rect 35 585 52 587
rect 72 585 75 587
rect 2 577 5 579
rect 35 577 52 579
rect 72 577 75 579
rect 2 569 5 571
rect 35 569 52 571
rect 72 569 75 571
rect 4 511 17 513
rect 37 511 51 513
rect 71 511 76 513
rect 4 503 17 505
rect 37 503 51 505
rect 71 503 76 505
rect 7 415 12 417
rect 52 415 64 417
rect 84 415 87 417
rect 7 407 12 409
rect 52 407 64 409
rect 84 407 87 409
rect 7 399 12 401
rect 52 399 64 401
rect 84 399 87 401
rect 7 391 12 393
rect 52 391 64 393
rect 84 391 87 393
rect 313 334 318 336
rect 358 334 370 336
rect 390 334 393 336
rect 4 330 7 332
rect 37 330 54 332
rect 74 330 77 332
rect 313 326 318 328
rect 358 326 370 328
rect 390 326 393 328
rect 4 322 7 324
rect 37 322 54 324
rect 74 322 77 324
rect 4 314 7 316
rect 37 314 54 316
rect 74 314 77 316
rect 313 318 318 320
rect 358 318 370 320
rect 390 318 393 320
rect 313 310 318 312
rect 358 310 370 312
rect 390 310 393 312
rect 4 259 17 261
rect 37 259 51 261
rect 71 259 76 261
rect 4 251 17 253
rect 37 251 51 253
rect 71 251 76 253
rect 5 167 8 169
rect 38 167 55 169
rect 75 167 78 169
rect 5 159 8 161
rect 38 159 55 161
rect 75 159 78 161
rect 5 151 8 153
rect 38 151 55 153
rect 75 151 78 153
rect 322 152 325 154
rect 355 152 372 154
rect 392 152 395 154
rect 322 144 325 146
rect 355 144 372 146
rect 392 144 395 146
rect 322 136 325 138
rect 355 136 372 138
rect 392 136 395 138
rect 5 96 18 98
rect 38 96 52 98
rect 72 96 77 98
rect 5 88 18 90
rect 38 88 52 90
rect 72 88 77 90
rect 3 13 16 15
rect 36 13 50 15
rect 70 13 75 15
rect 319 12 332 14
rect 352 12 366 14
rect 386 12 391 14
rect 3 5 16 7
rect 36 5 50 7
rect 70 5 75 7
rect 319 4 332 6
rect 352 4 366 6
rect 386 4 391 6
<< polycontact >>
rect 5 774 9 778
rect 5 766 9 770
rect 5 758 9 762
rect 5 750 9 754
rect 5 742 9 746
rect 1 679 5 683
rect 1 671 5 675
rect 1 663 5 667
rect 1 655 5 659
rect 300 635 304 639
rect 300 627 304 631
rect 300 619 304 623
rect 300 611 304 615
rect 300 603 304 607
rect -2 584 2 588
rect -2 576 2 580
rect -2 568 2 572
rect 0 510 4 514
rect 0 502 4 506
rect 3 414 7 418
rect 3 406 7 410
rect 3 398 7 402
rect 3 390 7 394
rect 0 329 4 333
rect 309 333 313 337
rect 0 321 4 325
rect 309 325 313 329
rect 0 313 4 317
rect 309 317 313 321
rect 309 309 313 313
rect 0 258 4 262
rect 0 250 4 254
rect 1 166 5 170
rect 1 158 5 162
rect 1 150 5 154
rect 318 151 322 155
rect 318 143 322 147
rect 318 135 322 139
rect 1 95 5 99
rect 1 87 5 91
rect -1 12 3 16
rect -1 4 3 8
rect 315 11 319 15
rect 315 3 319 7
<< metal1 >>
rect -409 845 258 850
rect 129 833 134 845
rect 68 805 233 810
rect 70 797 74 805
rect -418 779 -268 780
rect -418 776 5 779
rect 67 778 69 782
rect 101 778 103 782
rect -272 774 5 776
rect -272 683 -268 774
rect -248 766 5 771
rect 80 770 81 774
rect -227 758 5 763
rect 101 762 103 766
rect -182 753 5 754
rect -209 749 5 753
rect 80 754 81 758
rect -209 745 -144 749
rect 101 746 103 750
rect -9 741 5 746
rect 12 738 17 742
rect 12 727 16 738
rect 80 738 81 742
rect 12 723 152 727
rect 53 697 214 702
rect 53 687 57 697
rect 50 683 57 687
rect 82 683 129 687
rect -272 679 1 683
rect 53 679 57 683
rect -272 587 -268 679
rect 53 675 62 679
rect -2 674 1 675
rect -227 671 1 674
rect -2 666 1 667
rect -209 663 1 666
rect 53 663 57 675
rect 88 671 92 683
rect 82 667 92 671
rect 53 659 62 663
rect -9 656 1 659
rect -2 655 1 656
rect 88 655 92 667
rect 8 651 10 655
rect 82 651 92 655
rect 8 643 11 651
rect 8 640 153 643
rect 209 632 214 697
rect 228 640 233 805
rect 228 635 300 640
rect 362 639 364 643
rect 396 639 398 643
rect 209 627 300 632
rect 375 631 376 635
rect 167 620 300 624
rect 396 623 398 627
rect 46 619 300 620
rect 46 617 173 619
rect 201 610 300 615
rect 375 615 376 619
rect 35 588 41 592
rect 72 588 81 592
rect 201 590 206 610
rect 396 607 398 611
rect -272 584 -2 587
rect 41 584 45 588
rect -272 514 -268 584
rect 41 580 52 584
rect -226 576 -2 579
rect -148 568 -2 571
rect 43 568 47 580
rect 77 576 81 588
rect 72 572 81 576
rect 77 570 81 572
rect 43 564 52 568
rect 77 566 130 570
rect 16 554 20 564
rect 16 550 151 554
rect 8 526 130 530
rect 8 518 12 526
rect 71 519 151 523
rect 8 514 17 518
rect 71 514 75 519
rect -272 510 0 514
rect -191 503 -183 504
rect -176 503 0 506
rect -191 502 0 503
rect 8 502 12 514
rect 37 506 47 510
rect 43 502 47 506
rect -191 499 -172 502
rect -191 496 -183 499
rect 8 498 17 502
rect 43 498 51 502
rect 43 494 47 498
rect 202 494 206 590
rect 43 490 206 494
rect 219 602 300 607
rect 463 609 555 613
rect 219 486 224 602
rect 307 599 312 603
rect 307 591 311 599
rect 375 599 376 603
rect -406 478 224 486
rect 55 432 273 436
rect 55 422 59 432
rect 52 418 59 422
rect 84 418 130 422
rect -175 415 3 418
rect -408 414 3 415
rect 55 414 59 418
rect -408 409 -285 414
rect -280 410 -164 414
rect 55 410 64 414
rect -280 409 -184 410
rect -175 409 -164 410
rect -228 398 -177 401
rect -180 389 -176 390
rect -212 386 -176 389
rect -170 332 -164 409
rect -140 407 3 410
rect -140 404 -137 407
rect 0 406 3 407
rect -156 401 -137 404
rect -130 399 3 402
rect -130 393 -127 399
rect 0 398 3 399
rect 55 398 59 410
rect 90 406 94 418
rect 84 402 94 406
rect -156 390 -127 393
rect 55 394 64 398
rect -14 391 3 394
rect 0 390 3 391
rect 90 390 94 402
rect 10 386 12 390
rect 84 386 94 390
rect 10 375 13 386
rect 10 372 152 375
rect 108 345 216 348
rect 37 333 43 337
rect 74 333 83 337
rect -170 329 0 332
rect 43 329 47 333
rect -228 323 -180 326
rect -170 262 -164 329
rect 43 325 54 329
rect -156 321 0 324
rect -4 313 0 316
rect 45 313 49 325
rect 79 321 83 333
rect 213 328 216 345
rect 269 337 273 432
rect 361 355 436 359
rect 361 341 365 355
rect 358 337 365 341
rect 390 337 408 341
rect 269 333 309 337
rect 361 333 365 337
rect 361 329 370 333
rect 306 328 309 329
rect 213 325 309 328
rect 74 317 83 321
rect 306 320 309 321
rect 79 313 128 317
rect 182 317 309 320
rect 361 317 365 329
rect 396 325 400 337
rect 390 321 400 325
rect 45 309 54 313
rect 79 311 83 313
rect 18 302 22 309
rect 18 298 151 302
rect 8 274 130 278
rect 8 266 12 274
rect 71 270 75 271
rect 71 266 151 270
rect 8 262 17 266
rect 71 262 75 266
rect -170 258 0 262
rect -146 247 -7 251
rect -4 247 0 254
rect 8 250 12 262
rect 37 254 47 258
rect 43 250 47 254
rect -146 243 0 247
rect 8 246 17 250
rect 43 246 51 250
rect 43 236 47 246
rect 182 236 185 317
rect 361 313 370 317
rect 306 312 309 313
rect 273 309 309 312
rect 396 309 400 321
rect 43 232 188 236
rect 273 225 276 309
rect 316 305 318 309
rect 390 305 400 309
rect 316 301 319 305
rect 404 286 408 337
rect 432 316 436 355
rect 432 312 555 316
rect -402 217 -199 225
rect -191 217 280 225
rect 107 184 285 187
rect 38 170 44 174
rect 75 170 84 174
rect -404 164 -232 169
rect -227 166 1 169
rect 44 166 48 170
rect -227 164 -58 166
rect -136 99 -132 164
rect 44 162 55 166
rect -126 158 1 161
rect -126 139 -123 158
rect -14 150 1 153
rect 46 150 50 162
rect 80 158 84 170
rect 75 154 84 158
rect 80 152 84 154
rect 281 154 285 184
rect 355 155 361 159
rect 392 155 401 159
rect 46 146 55 150
rect 80 148 129 152
rect 281 151 318 154
rect 361 151 365 155
rect 361 147 372 151
rect 167 146 171 147
rect 19 137 23 146
rect 166 143 318 146
rect 19 133 150 137
rect 9 111 130 115
rect 9 103 13 111
rect 72 104 151 108
rect 9 99 18 103
rect 72 99 76 104
rect -136 95 1 99
rect -5 87 1 91
rect 9 87 13 99
rect 38 91 48 95
rect 44 87 48 91
rect 9 83 18 87
rect 44 83 52 87
rect 44 80 48 83
rect 167 80 171 143
rect 44 76 171 80
rect 295 135 318 138
rect 363 135 367 147
rect 397 143 401 155
rect 392 139 401 143
rect 429 141 553 144
rect 295 68 298 135
rect 363 131 372 135
rect 336 126 340 131
rect 397 116 401 139
rect -402 60 -154 68
rect -146 60 302 68
rect 295 59 298 60
rect 7 29 130 33
rect 156 32 186 36
rect 7 20 11 29
rect 182 28 390 32
rect 70 24 74 25
rect 70 20 152 24
rect 217 21 327 25
rect 7 16 16 20
rect 70 16 74 20
rect -401 5 -217 13
rect -209 11 -159 13
rect -154 12 -1 16
rect -154 11 -150 12
rect -209 7 -150 11
rect -209 5 -159 7
rect -21 4 -1 8
rect 7 4 11 16
rect 217 16 221 21
rect 323 19 327 21
rect 134 12 221 16
rect 268 13 315 17
rect 323 15 332 19
rect 386 15 390 28
rect 36 8 46 12
rect 42 4 46 8
rect -21 -27 -17 4
rect 7 0 16 4
rect 42 0 50 4
rect 42 -7 46 0
rect 268 -7 272 13
rect 311 11 315 13
rect 42 -11 272 -7
rect 295 3 315 7
rect 323 3 327 15
rect 352 7 362 11
rect 400 7 547 11
rect 358 3 362 7
rect 295 -27 299 3
rect 323 -1 332 3
rect 358 -1 366 3
rect 358 -7 362 -1
rect 400 -7 404 7
rect 358 -11 404 -7
rect -400 -28 300 -27
rect -400 -33 -161 -28
rect -156 -33 300 -28
rect -400 -35 300 -33
rect -403 -69 -159 -67
rect -21 -69 -17 -35
rect -403 -73 548 -69
rect -403 -75 -159 -73
rect -110 -74 -106 -73
rect 150 -166 156 -148
rect -431 -172 237 -166
<< m2contact >>
rect 129 828 134 833
rect 70 792 75 797
rect 69 778 74 783
rect 103 777 108 782
rect -253 766 -248 771
rect 75 769 80 774
rect -232 758 -227 763
rect 103 761 108 766
rect -217 745 -209 753
rect 75 753 80 758
rect -14 741 -9 746
rect 103 745 108 750
rect 75 737 80 742
rect 152 723 157 728
rect 129 683 134 688
rect -232 671 -227 676
rect -214 663 -209 668
rect -14 655 -9 660
rect 153 640 158 645
rect 364 639 369 644
rect 398 638 403 643
rect 370 630 375 635
rect 41 616 46 621
rect 398 622 403 627
rect 370 614 375 619
rect 41 588 46 593
rect -231 576 -226 581
rect -153 568 -148 573
rect 130 566 135 571
rect 151 550 156 555
rect 130 526 135 531
rect 151 519 156 524
rect -199 496 -191 504
rect 398 606 403 611
rect 458 609 463 614
rect 370 598 375 603
rect 307 586 312 591
rect 130 418 135 423
rect -285 409 -280 414
rect -233 398 -228 403
rect -182 401 -177 406
rect -217 386 -212 391
rect -161 400 -156 405
rect -161 390 -156 395
rect -19 391 -14 396
rect 152 372 157 377
rect 103 344 108 349
rect 43 333 48 338
rect -233 323 -228 328
rect -180 322 -175 327
rect -161 320 -156 325
rect -9 313 -4 318
rect 151 298 156 303
rect 130 274 135 279
rect 151 266 156 271
rect -154 243 -146 251
rect 316 296 321 301
rect 404 281 409 286
rect -199 217 -191 225
rect 102 183 107 188
rect 44 170 49 175
rect -232 164 -227 169
rect -19 150 -14 155
rect 361 155 366 160
rect 129 148 134 153
rect -127 134 -122 139
rect 130 111 135 116
rect 151 104 156 109
rect -10 87 -5 92
rect 424 140 429 145
rect 336 121 341 126
rect 397 111 402 116
rect -154 60 -146 68
rect 130 29 135 34
rect 151 32 156 37
rect 152 20 157 25
rect -217 5 -209 13
rect 129 12 134 17
rect -161 -33 -156 -28
rect -110 -69 -105 -64
rect 150 -148 156 -142
<< pdm12contact >>
rect -180 390 -175 395
rect 128 313 133 318
rect 150 133 155 138
<< metal2 >>
rect 70 783 74 792
rect 129 782 134 828
rect 70 774 74 778
rect 108 778 134 782
rect -285 766 -253 771
rect 70 770 75 774
rect -285 414 -280 766
rect -232 676 -227 758
rect 75 758 79 769
rect 103 766 107 777
rect -232 581 -227 671
rect -217 668 -209 745
rect -28 741 -14 746
rect 75 742 79 753
rect 103 750 107 761
rect -217 663 -214 668
rect -232 576 -231 581
rect -232 403 -227 576
rect -228 398 -227 403
rect -232 328 -227 398
rect -228 323 -227 328
rect -232 169 -227 323
rect -217 391 -209 663
rect 129 688 134 778
rect -117 659 -14 660
rect -118 657 -14 659
rect -212 386 -209 391
rect -217 145 -209 386
rect -199 225 -191 496
rect -177 402 -161 405
rect -175 391 -161 394
rect -175 322 -161 325
rect -152 251 -149 568
rect -118 317 -114 657
rect 41 596 44 616
rect 40 593 44 596
rect 129 582 134 683
rect 150 728 156 794
rect 150 723 152 728
rect 150 645 156 723
rect 365 658 462 662
rect 150 640 153 645
rect 365 644 369 658
rect 150 590 156 640
rect 365 635 369 639
rect 403 639 412 643
rect 365 631 370 635
rect 370 619 374 630
rect 398 627 402 638
rect 370 603 374 614
rect 398 611 402 622
rect 150 586 307 590
rect 129 579 144 582
rect 129 578 140 579
rect 129 571 134 578
rect 129 566 130 571
rect 129 531 134 566
rect 150 555 156 586
rect 408 578 412 639
rect 458 614 462 658
rect 254 574 412 578
rect 150 550 151 555
rect 129 526 130 531
rect 129 423 134 526
rect 150 524 156 550
rect 150 519 151 524
rect 129 418 130 423
rect -23 392 -19 395
rect 43 344 103 347
rect 43 341 46 344
rect 42 338 46 341
rect 129 318 134 418
rect -118 314 -9 317
rect -172 147 -171 149
rect -154 151 -146 243
rect -166 148 -129 151
rect -172 145 -166 147
rect -218 142 -166 145
rect -217 139 -166 142
rect -217 13 -209 139
rect -154 68 -146 148
rect -128 139 -125 147
rect -128 135 -127 139
rect -118 91 -114 314
rect 133 313 134 318
rect 129 289 134 313
rect 150 377 156 519
rect 150 372 152 377
rect 150 303 156 372
rect 150 298 151 303
rect 156 298 316 300
rect 150 297 316 298
rect 129 286 143 289
rect 129 285 139 286
rect 129 279 134 285
rect 129 274 130 279
rect 44 183 102 186
rect 44 178 47 183
rect 43 175 47 178
rect -23 151 -19 154
rect 129 153 134 274
rect 129 116 134 148
rect 150 271 156 297
rect 210 281 404 285
rect 150 266 151 271
rect 150 138 156 266
rect 360 172 427 175
rect 360 163 363 172
rect 360 160 364 163
rect 424 145 427 172
rect 155 133 156 138
rect 150 125 156 133
rect 150 121 336 125
rect 129 111 130 116
rect 135 111 140 115
rect -133 87 -10 91
rect -133 -29 -129 87
rect 129 34 134 111
rect 150 109 156 121
rect 234 111 397 115
rect 150 104 151 109
rect 150 37 156 104
rect 129 29 130 34
rect 150 32 151 37
rect 129 17 134 29
rect 129 -16 134 12
rect 150 25 156 32
rect 150 20 152 25
rect -156 -33 -129 -29
rect -110 -64 -106 -57
rect 150 -142 156 20
<< m3contact >>
rect -33 741 -28 746
rect 140 574 145 579
rect 249 574 254 579
rect -28 391 -23 396
rect -171 147 -166 152
rect -129 147 -124 152
rect 139 281 144 286
rect -28 150 -23 155
rect 205 281 210 286
rect 140 111 145 116
rect 229 111 234 116
rect -110 -57 -105 -52
<< metal3 >>
rect -34 746 -27 747
rect -110 741 -33 746
rect -28 741 -27 746
rect -109 395 -105 741
rect -34 740 -27 741
rect 139 579 146 580
rect 139 574 140 579
rect 145 578 146 579
rect 248 579 255 580
rect 248 578 249 579
rect 145 574 249 578
rect 254 574 255 579
rect 139 573 146 574
rect 248 573 255 574
rect -29 396 -22 397
rect -29 395 -28 396
rect -109 392 -28 395
rect -109 154 -105 392
rect -29 391 -28 392
rect -23 391 -22 396
rect -29 390 -22 391
rect 138 286 145 287
rect 138 281 139 286
rect 144 285 145 286
rect 204 286 211 287
rect 204 285 205 286
rect 144 281 205 285
rect 210 281 211 286
rect 138 280 145 281
rect 204 280 211 281
rect -29 155 -22 156
rect -29 154 -28 155
rect -172 152 -165 153
rect -172 147 -171 152
rect -166 151 -165 152
rect -130 152 -123 153
rect -130 151 -129 152
rect -166 148 -129 151
rect -166 147 -165 148
rect -172 146 -165 147
rect -130 147 -129 148
rect -124 147 -123 152
rect -130 146 -123 147
rect -109 151 -28 154
rect -109 -51 -105 151
rect -29 150 -28 151
rect -23 150 -22 155
rect -29 149 -22 150
rect 139 116 146 117
rect 139 111 140 116
rect 145 115 146 116
rect 228 116 235 117
rect 228 115 229 116
rect 145 111 229 115
rect 234 111 235 116
rect 139 110 146 111
rect 228 110 235 111
rect -111 -52 -104 -51
rect -111 -57 -110 -52
rect -105 -57 -104 -52
rect -111 -58 -104 -57
<< labels >>
rlabel space -407 -88 -388 -62 1 G0
rlabel space -403 -45 -384 -19 1 G1
rlabel space -403 -1 -384 25 1 P1
rlabel space -404 49 -385 75 1 G2
rlabel space -410 155 -391 181 1 P2
rlabel space -404 205 -385 231 1 G3
rlabel space -412 397 -393 423 1 P3
rlabel space -409 466 -390 492 1 G4
rlabel space -423 766 -404 792 1 P4
rlabel space 528 -86 557 -60 1 C1
rlabel space 527 -4 556 22 1 C2
rlabel space 535 128 564 154 1 C3
rlabel space 536 301 565 327 1 C4
rlabel space 535 597 564 623 1 C5
rlabel space -433 -180 -404 -154 1 ground
rlabel space -412 835 -383 861 5 power
<< end >>
