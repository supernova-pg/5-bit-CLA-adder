magic
tech scmos
timestamp 1764703505
<< nwell >>
rect 1 28 62 60
rect 91 7 123 39
rect 135 33 160 65
rect 217 28 278 60
rect 307 7 339 39
rect 351 33 376 65
rect 433 28 494 60
rect 523 7 555 39
rect 567 33 592 65
rect 649 28 710 60
rect 739 7 771 39
rect 783 33 808 65
rect 865 28 926 60
rect 955 7 987 39
rect 999 33 1024 65
<< ntransistor >>
rect 102 47 104 67
rect 110 47 112 67
rect 12 12 14 22
rect 40 11 42 21
rect 49 11 51 21
rect 318 47 320 67
rect 326 47 328 67
rect 146 17 148 27
rect 228 12 230 22
rect 256 11 258 21
rect 265 11 267 21
rect 534 47 536 67
rect 542 47 544 67
rect 362 17 364 27
rect 444 12 446 22
rect 472 11 474 21
rect 481 11 483 21
rect 750 47 752 67
rect 758 47 760 67
rect 578 17 580 27
rect 660 12 662 22
rect 688 11 690 21
rect 697 11 699 21
rect 966 47 968 67
rect 974 47 976 67
rect 794 17 796 27
rect 876 12 878 22
rect 904 11 906 21
rect 913 11 915 21
rect 1010 17 1012 27
<< ptransistor >>
rect 12 34 14 54
rect 40 34 42 54
rect 49 34 51 54
rect 146 39 148 59
rect 102 13 104 33
rect 110 13 112 33
rect 228 34 230 54
rect 256 34 258 54
rect 265 34 267 54
rect 362 39 364 59
rect 318 13 320 33
rect 326 13 328 33
rect 444 34 446 54
rect 472 34 474 54
rect 481 34 483 54
rect 578 39 580 59
rect 534 13 536 33
rect 542 13 544 33
rect 660 34 662 54
rect 688 34 690 54
rect 697 34 699 54
rect 794 39 796 59
rect 750 13 752 33
rect 758 13 760 33
rect 876 34 878 54
rect 904 34 906 54
rect 913 34 915 54
rect 1010 39 1012 59
rect 966 13 968 33
rect 974 13 976 33
<< ndiffusion >>
rect 101 47 102 67
rect 104 47 105 67
rect 109 47 110 67
rect 112 47 113 67
rect 7 16 12 22
rect 11 12 12 16
rect 14 16 19 22
rect 14 12 15 16
rect 35 15 40 21
rect 39 11 40 15
rect 42 17 43 21
rect 47 17 49 21
rect 42 11 49 17
rect 51 17 52 21
rect 51 11 56 17
rect 317 47 318 67
rect 320 47 321 67
rect 325 47 326 67
rect 328 47 329 67
rect 141 21 146 27
rect 145 17 146 21
rect 148 23 149 27
rect 148 17 153 23
rect 223 16 228 22
rect 227 12 228 16
rect 230 16 235 22
rect 230 12 231 16
rect 251 15 256 21
rect 255 11 256 15
rect 258 17 259 21
rect 263 17 265 21
rect 258 11 265 17
rect 267 17 268 21
rect 267 11 272 17
rect 533 47 534 67
rect 536 47 537 67
rect 541 47 542 67
rect 544 47 545 67
rect 357 21 362 27
rect 361 17 362 21
rect 364 23 365 27
rect 364 17 369 23
rect 439 16 444 22
rect 443 12 444 16
rect 446 16 451 22
rect 446 12 447 16
rect 467 15 472 21
rect 471 11 472 15
rect 474 17 475 21
rect 479 17 481 21
rect 474 11 481 17
rect 483 17 484 21
rect 483 11 488 17
rect 749 47 750 67
rect 752 47 753 67
rect 757 47 758 67
rect 760 47 761 67
rect 573 21 578 27
rect 577 17 578 21
rect 580 23 581 27
rect 580 17 585 23
rect 655 16 660 22
rect 659 12 660 16
rect 662 16 667 22
rect 662 12 663 16
rect 683 15 688 21
rect 687 11 688 15
rect 690 17 691 21
rect 695 17 697 21
rect 690 11 697 17
rect 699 17 700 21
rect 699 11 704 17
rect 965 47 966 67
rect 968 47 969 67
rect 973 47 974 67
rect 976 47 977 67
rect 789 21 794 27
rect 793 17 794 21
rect 796 23 797 27
rect 796 17 801 23
rect 871 16 876 22
rect 875 12 876 16
rect 878 16 883 22
rect 878 12 879 16
rect 899 15 904 21
rect 903 11 904 15
rect 906 17 907 21
rect 911 17 913 21
rect 906 11 913 17
rect 915 17 916 21
rect 915 11 920 17
rect 1005 21 1010 27
rect 1009 17 1010 21
rect 1012 23 1013 27
rect 1012 17 1017 23
<< pdiffusion >>
rect 7 38 12 54
rect 11 34 12 38
rect 14 50 15 54
rect 14 34 19 50
rect 39 50 40 54
rect 35 34 40 50
rect 42 40 49 54
rect 42 36 43 40
rect 47 36 49 40
rect 42 34 49 36
rect 51 38 56 54
rect 145 55 146 59
rect 51 34 52 38
rect 141 39 146 55
rect 148 43 153 59
rect 148 39 149 43
rect 101 13 102 33
rect 104 13 105 33
rect 109 13 110 33
rect 112 13 113 33
rect 223 38 228 54
rect 227 34 228 38
rect 230 50 231 54
rect 230 34 235 50
rect 255 50 256 54
rect 251 34 256 50
rect 258 40 265 54
rect 258 36 259 40
rect 263 36 265 40
rect 258 34 265 36
rect 267 38 272 54
rect 361 55 362 59
rect 267 34 268 38
rect 357 39 362 55
rect 364 43 369 59
rect 364 39 365 43
rect 317 13 318 33
rect 320 13 321 33
rect 325 13 326 33
rect 328 13 329 33
rect 439 38 444 54
rect 443 34 444 38
rect 446 50 447 54
rect 446 34 451 50
rect 471 50 472 54
rect 467 34 472 50
rect 474 40 481 54
rect 474 36 475 40
rect 479 36 481 40
rect 474 34 481 36
rect 483 38 488 54
rect 577 55 578 59
rect 483 34 484 38
rect 573 39 578 55
rect 580 43 585 59
rect 580 39 581 43
rect 533 13 534 33
rect 536 13 537 33
rect 541 13 542 33
rect 544 13 545 33
rect 655 38 660 54
rect 659 34 660 38
rect 662 50 663 54
rect 662 34 667 50
rect 687 50 688 54
rect 683 34 688 50
rect 690 40 697 54
rect 690 36 691 40
rect 695 36 697 40
rect 690 34 697 36
rect 699 38 704 54
rect 793 55 794 59
rect 699 34 700 38
rect 789 39 794 55
rect 796 43 801 59
rect 796 39 797 43
rect 749 13 750 33
rect 752 13 753 33
rect 757 13 758 33
rect 760 13 761 33
rect 871 38 876 54
rect 875 34 876 38
rect 878 50 879 54
rect 878 34 883 50
rect 903 50 904 54
rect 899 34 904 50
rect 906 40 913 54
rect 906 36 907 40
rect 911 36 913 40
rect 906 34 913 36
rect 915 38 920 54
rect 1009 55 1010 59
rect 915 34 916 38
rect 1005 39 1010 55
rect 1012 43 1017 59
rect 1012 39 1013 43
rect 965 13 966 33
rect 968 13 969 33
rect 973 13 974 33
rect 976 13 977 33
<< ndcontact >>
rect 97 47 101 67
rect 105 47 109 67
rect 113 47 117 67
rect 7 12 11 16
rect 15 12 19 16
rect 35 11 39 15
rect 43 17 47 21
rect 52 17 56 21
rect 313 47 317 67
rect 321 47 325 67
rect 329 47 333 67
rect 141 17 145 21
rect 149 23 153 27
rect 223 12 227 16
rect 231 12 235 16
rect 251 11 255 15
rect 259 17 263 21
rect 268 17 272 21
rect 529 47 533 67
rect 537 47 541 67
rect 545 47 549 67
rect 357 17 361 21
rect 365 23 369 27
rect 439 12 443 16
rect 447 12 451 16
rect 467 11 471 15
rect 475 17 479 21
rect 484 17 488 21
rect 745 47 749 67
rect 753 47 757 67
rect 761 47 765 67
rect 573 17 577 21
rect 581 23 585 27
rect 655 12 659 16
rect 663 12 667 16
rect 683 11 687 15
rect 691 17 695 21
rect 700 17 704 21
rect 961 47 965 67
rect 969 47 973 67
rect 977 47 981 67
rect 789 17 793 21
rect 797 23 801 27
rect 871 12 875 16
rect 879 12 883 16
rect 899 11 903 15
rect 907 17 911 21
rect 916 17 920 21
rect 1005 17 1009 21
rect 1013 23 1017 27
<< pdcontact >>
rect 7 34 11 38
rect 15 50 19 54
rect 35 50 39 54
rect 43 36 47 40
rect 141 55 145 59
rect 52 34 56 38
rect 149 39 153 43
rect 97 13 101 33
rect 105 13 109 33
rect 113 13 117 33
rect 223 34 227 38
rect 231 50 235 54
rect 251 50 255 54
rect 259 36 263 40
rect 357 55 361 59
rect 268 34 272 38
rect 365 39 369 43
rect 313 13 317 33
rect 321 13 325 33
rect 329 13 333 33
rect 439 34 443 38
rect 447 50 451 54
rect 467 50 471 54
rect 475 36 479 40
rect 573 55 577 59
rect 484 34 488 38
rect 581 39 585 43
rect 529 13 533 33
rect 537 13 541 33
rect 545 13 549 33
rect 655 34 659 38
rect 663 50 667 54
rect 683 50 687 54
rect 691 36 695 40
rect 789 55 793 59
rect 700 34 704 38
rect 797 39 801 43
rect 745 13 749 33
rect 753 13 757 33
rect 761 13 765 33
rect 871 34 875 38
rect 879 50 883 54
rect 899 50 903 54
rect 907 36 911 40
rect 1005 55 1009 59
rect 916 34 920 38
rect 1013 39 1017 43
rect 961 13 965 33
rect 969 13 973 33
rect 977 13 981 33
<< polysilicon >>
rect 102 67 104 72
rect 110 67 112 72
rect 318 67 320 72
rect 326 67 328 72
rect 534 67 536 72
rect 542 67 544 72
rect 750 67 752 72
rect 758 67 760 72
rect 966 67 968 72
rect 974 67 976 72
rect 12 54 14 58
rect 40 54 42 57
rect 49 54 51 66
rect 146 59 148 63
rect 12 22 14 34
rect 40 21 42 34
rect 49 28 51 34
rect 102 33 104 47
rect 110 33 112 47
rect 228 54 230 58
rect 256 54 258 57
rect 265 54 267 66
rect 49 21 51 25
rect 12 8 14 12
rect 146 27 148 39
rect 362 59 364 63
rect 228 22 230 34
rect 146 13 148 17
rect 40 8 42 11
rect 49 9 51 11
rect 50 5 51 9
rect 49 4 51 5
rect 102 0 104 13
rect 110 0 112 13
rect 256 21 258 34
rect 265 28 267 34
rect 318 33 320 47
rect 326 33 328 47
rect 444 54 446 58
rect 472 54 474 57
rect 481 54 483 66
rect 265 21 267 25
rect 228 8 230 12
rect 362 27 364 39
rect 578 59 580 63
rect 444 22 446 34
rect 362 13 364 17
rect 256 8 258 11
rect 265 9 267 11
rect 266 5 267 9
rect 265 4 267 5
rect 318 0 320 13
rect 326 0 328 13
rect 472 21 474 34
rect 481 28 483 34
rect 534 33 536 47
rect 542 33 544 47
rect 660 54 662 58
rect 688 54 690 57
rect 697 54 699 66
rect 481 21 483 25
rect 444 8 446 12
rect 578 27 580 39
rect 794 59 796 63
rect 660 22 662 34
rect 578 13 580 17
rect 472 8 474 11
rect 481 9 483 11
rect 482 5 483 9
rect 481 4 483 5
rect 534 0 536 13
rect 542 0 544 13
rect 688 21 690 34
rect 697 28 699 34
rect 750 33 752 47
rect 758 33 760 47
rect 876 54 878 58
rect 904 54 906 57
rect 913 54 915 66
rect 697 21 699 25
rect 660 8 662 12
rect 794 27 796 39
rect 1010 59 1012 63
rect 876 22 878 34
rect 794 13 796 17
rect 688 8 690 11
rect 697 9 699 11
rect 698 5 699 9
rect 697 4 699 5
rect 750 0 752 13
rect 758 0 760 13
rect 904 21 906 34
rect 913 28 915 34
rect 966 33 968 47
rect 974 33 976 47
rect 913 21 915 25
rect 876 8 878 12
rect 1010 27 1012 39
rect 1010 13 1012 17
rect 904 8 906 11
rect 913 9 915 11
rect 914 5 915 9
rect 913 4 915 5
rect 966 0 968 13
rect 974 0 976 13
<< polycontact >>
rect 45 61 49 65
rect 261 61 265 65
rect 14 23 18 27
rect 36 23 40 27
rect 142 28 146 32
rect 477 61 481 65
rect 230 23 234 27
rect 252 23 256 27
rect 46 5 50 9
rect 358 28 362 32
rect 693 61 697 65
rect 446 23 450 27
rect 468 23 472 27
rect 262 5 266 9
rect 574 28 578 32
rect 909 61 913 65
rect 662 23 666 27
rect 684 23 688 27
rect 478 5 482 9
rect 790 28 794 32
rect 878 23 882 27
rect 900 23 904 27
rect 694 5 698 9
rect 1006 28 1010 32
rect 910 5 914 9
rect 101 -4 105 0
rect 109 -4 113 0
rect 317 -4 321 0
rect 325 -4 329 0
rect 533 -4 537 0
rect 541 -4 545 0
rect 749 -4 753 0
rect 757 -4 761 0
rect 965 -4 969 0
rect 973 -4 977 0
<< metal1 >>
rect 31 74 34 95
rect 101 86 104 94
rect 101 83 167 86
rect 79 67 101 71
rect 131 67 154 69
rect 0 63 14 66
rect 15 54 19 61
rect 30 61 45 64
rect 30 54 33 61
rect 22 51 35 54
rect 7 18 10 34
rect 22 27 25 51
rect 44 33 47 36
rect 18 24 25 27
rect 6 16 10 18
rect 6 13 7 16
rect 0 4 15 7
rect 9 -14 12 4
rect 22 -11 25 24
rect 33 23 36 26
rect 44 21 47 28
rect 52 27 55 34
rect 79 29 82 67
rect 136 66 154 67
rect 141 59 144 66
rect 159 66 160 69
rect 113 43 117 47
rect 105 39 131 43
rect 105 33 109 39
rect 52 25 70 27
rect 52 24 59 25
rect 52 21 55 24
rect 64 24 70 25
rect 29 10 35 14
rect 34 8 35 10
rect 34 5 46 8
rect 67 5 70 24
rect 127 32 131 39
rect 150 32 153 39
rect 164 32 167 83
rect 247 74 250 95
rect 317 86 320 94
rect 317 83 383 86
rect 218 66 221 74
rect 295 67 317 71
rect 347 67 370 69
rect 216 63 230 66
rect 231 54 235 61
rect 246 61 261 64
rect 246 54 249 61
rect 238 51 251 54
rect 127 29 142 32
rect 150 29 167 32
rect 150 27 153 29
rect 124 13 127 21
rect 97 8 101 13
rect 113 10 127 13
rect 223 18 226 34
rect 238 27 241 51
rect 260 33 263 36
rect 234 24 241 27
rect 141 12 144 17
rect 113 9 126 10
rect 134 9 157 12
rect 222 16 226 18
rect 222 13 223 16
rect 113 8 124 9
rect 60 2 70 5
rect 91 7 124 8
rect 91 4 122 7
rect 134 6 137 9
rect 60 1 63 2
rect 132 3 137 6
rect 216 4 231 7
rect 35 -2 63 1
rect 35 -10 38 -2
rect 101 -8 105 -4
rect 22 -14 29 -11
rect 35 -13 86 -10
rect 101 -10 104 -8
rect 91 -13 104 -10
rect 26 -20 29 -14
rect 109 -20 113 -4
rect 225 -14 228 4
rect 238 -11 241 24
rect 249 23 252 26
rect 260 21 263 28
rect 268 27 271 34
rect 295 29 298 67
rect 352 66 370 67
rect 357 59 360 66
rect 375 66 376 69
rect 329 43 333 47
rect 321 39 347 43
rect 321 33 325 39
rect 268 25 286 27
rect 268 24 275 25
rect 268 21 271 24
rect 280 24 286 25
rect 245 10 251 14
rect 250 8 251 10
rect 250 5 262 8
rect 283 5 286 24
rect 343 32 347 39
rect 366 32 369 39
rect 380 32 383 83
rect 463 74 466 95
rect 533 86 536 94
rect 533 83 599 86
rect 433 66 436 73
rect 511 67 533 71
rect 563 67 586 69
rect 432 63 446 66
rect 447 54 451 61
rect 462 61 477 64
rect 462 54 465 61
rect 454 51 467 54
rect 343 29 358 32
rect 366 29 383 32
rect 366 27 369 29
rect 340 13 343 21
rect 313 8 317 13
rect 329 10 343 13
rect 439 18 442 34
rect 454 27 457 51
rect 476 33 479 36
rect 450 24 457 27
rect 357 12 360 17
rect 438 16 442 18
rect 438 13 439 16
rect 329 9 342 10
rect 350 9 376 12
rect 329 8 340 9
rect 276 2 286 5
rect 307 7 340 8
rect 307 4 338 7
rect 350 6 353 9
rect 276 1 279 2
rect 348 3 353 6
rect 432 4 447 7
rect 251 -2 279 1
rect 251 -10 254 -2
rect 317 -8 321 -4
rect 238 -14 245 -11
rect 251 -13 302 -10
rect 317 -10 320 -8
rect 307 -13 320 -10
rect 26 -23 113 -20
rect 242 -20 245 -14
rect 325 -20 329 -4
rect 441 -14 444 4
rect 454 -11 457 24
rect 465 23 468 26
rect 476 21 479 28
rect 484 27 487 34
rect 511 29 514 67
rect 568 66 586 67
rect 573 59 576 66
rect 591 66 592 69
rect 545 43 549 47
rect 537 39 563 43
rect 537 33 541 39
rect 484 25 502 27
rect 484 24 491 25
rect 484 21 487 24
rect 496 24 502 25
rect 461 10 467 14
rect 466 8 467 10
rect 466 5 478 8
rect 499 5 502 24
rect 559 32 563 39
rect 582 32 585 39
rect 596 32 599 83
rect 679 74 682 95
rect 749 86 752 94
rect 749 83 815 86
rect 650 66 653 74
rect 727 67 749 71
rect 779 67 802 69
rect 648 63 662 66
rect 663 54 667 61
rect 678 61 693 64
rect 678 54 681 61
rect 670 51 683 54
rect 559 29 574 32
rect 582 29 599 32
rect 582 27 585 29
rect 556 13 559 21
rect 529 8 533 13
rect 545 10 559 13
rect 655 18 658 34
rect 670 27 673 51
rect 692 33 695 36
rect 666 24 673 27
rect 573 12 576 17
rect 654 16 658 18
rect 654 13 655 16
rect 545 9 558 10
rect 566 9 592 12
rect 545 8 556 9
rect 492 2 502 5
rect 523 7 556 8
rect 523 4 554 7
rect 566 6 569 9
rect 492 1 495 2
rect 564 3 569 6
rect 648 4 663 7
rect 467 -2 495 1
rect 467 -10 470 -2
rect 533 -8 537 -4
rect 454 -14 461 -11
rect 467 -13 518 -10
rect 533 -10 536 -8
rect 523 -13 536 -10
rect 242 -23 329 -20
rect 458 -20 461 -14
rect 541 -20 545 -4
rect 657 -14 660 4
rect 670 -11 673 24
rect 681 23 684 26
rect 692 21 695 28
rect 700 27 703 34
rect 727 29 730 67
rect 784 66 802 67
rect 789 59 792 66
rect 807 66 808 69
rect 761 43 765 47
rect 753 39 779 43
rect 753 33 757 39
rect 700 25 718 27
rect 700 24 707 25
rect 700 21 703 24
rect 712 24 718 25
rect 677 10 683 14
rect 682 8 683 10
rect 682 5 694 8
rect 715 5 718 24
rect 775 32 779 39
rect 798 32 801 39
rect 812 32 815 83
rect 895 74 898 95
rect 965 86 968 94
rect 965 83 1031 86
rect 867 66 870 74
rect 943 67 965 71
rect 995 67 1018 69
rect 864 63 878 66
rect 879 54 883 61
rect 894 61 909 64
rect 894 54 897 61
rect 886 51 899 54
rect 775 29 790 32
rect 798 29 815 32
rect 798 27 801 29
rect 772 13 775 21
rect 745 8 749 13
rect 761 10 775 13
rect 871 18 874 34
rect 886 27 889 51
rect 908 33 911 36
rect 882 24 889 27
rect 789 12 792 17
rect 870 16 874 18
rect 870 13 871 16
rect 761 9 774 10
rect 782 9 808 12
rect 761 8 772 9
rect 708 2 718 5
rect 739 7 772 8
rect 739 4 770 7
rect 782 6 785 9
rect 708 1 711 2
rect 780 3 785 6
rect 864 4 879 7
rect 683 -2 711 1
rect 683 -10 686 -2
rect 749 -8 753 -4
rect 670 -14 677 -11
rect 683 -13 734 -10
rect 749 -10 752 -8
rect 739 -13 752 -10
rect 458 -23 545 -20
rect 674 -20 677 -14
rect 757 -20 761 -4
rect 873 -14 876 4
rect 886 -11 889 24
rect 897 23 900 26
rect 908 21 911 28
rect 916 27 919 34
rect 943 29 946 67
rect 1000 66 1018 67
rect 1005 59 1008 66
rect 1023 66 1024 69
rect 977 43 981 47
rect 969 39 995 43
rect 969 33 973 39
rect 916 25 934 27
rect 916 24 923 25
rect 916 21 919 24
rect 928 24 934 25
rect 893 10 899 14
rect 898 8 899 10
rect 898 5 910 8
rect 931 5 934 24
rect 991 32 995 39
rect 1014 32 1017 39
rect 1028 32 1031 83
rect 991 29 1006 32
rect 1014 29 1031 32
rect 1014 27 1017 29
rect 988 13 991 21
rect 961 8 965 13
rect 977 10 991 13
rect 1005 12 1008 17
rect 977 9 990 10
rect 998 9 1024 12
rect 977 8 988 9
rect 924 2 934 5
rect 955 7 988 8
rect 955 4 986 7
rect 998 6 1001 9
rect 924 1 927 2
rect 996 3 1001 6
rect 899 -2 927 1
rect 899 -10 902 -2
rect 965 -8 969 -4
rect 886 -14 893 -11
rect 899 -13 950 -10
rect 965 -10 968 -8
rect 955 -13 968 -10
rect 674 -23 761 -20
rect 890 -20 893 -14
rect 973 -20 977 -4
rect 890 -23 977 -20
rect 109 -30 113 -23
rect 88 -54 91 -33
rect 100 -34 113 -30
rect 325 -30 329 -23
rect 100 -54 104 -34
rect 304 -52 307 -33
rect 316 -34 329 -30
rect 541 -30 545 -23
rect 316 -52 320 -34
rect 520 -52 523 -33
rect 532 -34 545 -30
rect 757 -30 761 -23
rect 532 -52 536 -34
rect 736 -49 739 -33
rect 748 -34 761 -30
rect 973 -30 977 -23
rect 748 -49 752 -34
rect 952 -50 955 -33
rect 964 -34 977 -30
rect 964 -50 968 -34
<< m2contact >>
rect 30 69 35 74
rect 14 61 19 66
rect 43 28 48 33
rect 1 13 6 18
rect 131 62 136 67
rect 154 65 159 70
rect 78 24 83 29
rect 29 5 34 10
rect 217 74 222 79
rect 246 69 251 74
rect 230 61 235 66
rect 123 21 128 26
rect 259 28 264 33
rect 157 9 162 14
rect 217 13 222 18
rect 127 1 132 6
rect 86 -13 91 -8
rect 9 -19 14 -14
rect 347 62 352 67
rect 370 65 375 70
rect 294 24 299 29
rect 245 5 250 10
rect 432 73 437 78
rect 462 69 467 74
rect 446 61 451 66
rect 339 21 344 26
rect 475 28 480 33
rect 433 13 438 18
rect 343 1 348 6
rect 302 -13 307 -8
rect 225 -19 230 -14
rect 563 62 568 67
rect 586 65 591 70
rect 510 24 515 29
rect 461 5 466 10
rect 649 74 654 79
rect 678 69 683 74
rect 662 61 667 66
rect 555 21 560 26
rect 691 28 696 33
rect 649 13 654 18
rect 559 1 564 6
rect 518 -13 523 -8
rect 441 -19 446 -14
rect 779 62 784 67
rect 802 65 807 70
rect 726 24 731 29
rect 677 5 682 10
rect 866 74 871 79
rect 894 69 899 74
rect 878 61 883 66
rect 771 21 776 26
rect 907 28 912 33
rect 865 13 870 18
rect 775 1 780 6
rect 734 -13 739 -8
rect 657 -19 662 -14
rect 995 62 1000 67
rect 1018 65 1023 70
rect 942 24 947 29
rect 893 5 898 10
rect 987 21 992 26
rect 991 1 996 6
rect 950 -13 955 -8
rect 873 -19 878 -14
rect 87 -33 92 -28
rect 303 -33 308 -28
rect 519 -33 524 -28
rect 735 -33 740 -28
rect 951 -33 956 -28
<< metal2 >>
rect 133 76 217 77
rect 127 74 217 76
rect 127 72 136 74
rect 35 69 69 72
rect 155 70 158 74
rect 19 62 20 66
rect 66 32 69 69
rect 349 76 432 77
rect 343 74 432 76
rect 343 72 352 74
rect 251 69 285 72
rect 371 70 374 74
rect 48 29 69 32
rect 78 19 81 24
rect 132 24 135 62
rect 235 62 236 66
rect 282 32 285 69
rect 565 76 649 77
rect 559 74 649 76
rect 559 72 568 74
rect 467 69 501 72
rect 587 70 590 74
rect 264 29 285 32
rect 128 21 135 24
rect 294 19 297 24
rect 348 24 351 62
rect 451 62 452 66
rect 498 32 501 69
rect 781 76 866 77
rect 775 74 866 76
rect 775 72 784 74
rect 683 69 717 72
rect 803 70 806 74
rect 480 29 501 32
rect 344 21 351 24
rect 510 19 513 24
rect 564 24 567 62
rect 667 62 668 66
rect 714 32 717 69
rect 997 76 1022 77
rect 991 74 1022 76
rect 991 72 1000 74
rect 899 69 933 72
rect 1019 70 1022 74
rect 696 29 717 32
rect 560 21 567 24
rect 726 19 729 24
rect 780 24 783 62
rect 883 62 884 66
rect 930 32 933 69
rect 912 29 933 32
rect 776 21 783 24
rect 942 19 945 24
rect 996 24 999 62
rect 992 21 999 24
rect 2 -5 5 13
rect 29 -5 32 5
rect 2 -8 32 -5
rect 10 -24 13 -19
rect 87 -28 90 -13
rect 158 -37 161 9
rect 218 -5 221 13
rect 245 -5 248 5
rect 218 -8 248 -5
rect 226 -24 229 -19
rect 303 -28 306 -13
rect 343 -37 346 1
rect 434 -5 437 13
rect 461 -5 464 5
rect 434 -8 464 -5
rect 442 -24 445 -19
rect 519 -28 522 -13
rect 560 -37 563 1
rect 650 -5 653 13
rect 677 -5 680 5
rect 650 -8 680 -5
rect 658 -24 661 -19
rect 735 -28 738 -13
rect 158 -38 563 -37
rect 776 -38 779 1
rect 866 -5 869 13
rect 893 -5 896 5
rect 866 -8 896 -5
rect 874 -24 877 -19
rect 951 -28 954 -13
rect 991 -38 994 1
rect 158 -40 994 -38
rect 560 -41 994 -40
rect 560 -44 563 -41
<< m3contact >>
rect 122 72 127 77
rect 20 62 25 67
rect 338 72 343 77
rect 236 62 241 67
rect 554 72 559 77
rect 452 62 457 67
rect 770 72 775 77
rect 668 62 673 67
rect 986 72 991 77
rect 884 62 889 67
rect 77 14 82 19
rect 127 6 132 11
rect 293 14 298 19
rect 509 14 514 19
rect 725 14 730 19
rect 941 14 946 19
rect 9 -29 14 -24
rect 343 6 348 11
rect 225 -29 230 -24
rect 559 6 564 11
rect 441 -29 446 -24
rect 775 6 780 11
rect 657 -29 662 -24
rect 991 6 996 11
rect 873 -29 878 -24
<< m123contact >>
rect 28 22 33 27
rect 59 20 64 25
rect 244 22 249 27
rect 275 20 280 25
rect 460 22 465 27
rect 491 20 496 25
rect 676 22 681 27
rect 707 20 712 25
rect 892 22 897 27
rect 923 20 928 25
<< metal3 >>
rect 121 77 128 78
rect 121 72 122 77
rect 127 72 128 77
rect 121 71 128 72
rect 337 77 344 78
rect 337 72 338 77
rect 343 72 344 77
rect 337 71 344 72
rect 553 77 560 78
rect 553 72 554 77
rect 559 72 560 77
rect 553 71 560 72
rect 769 77 776 78
rect 769 72 770 77
rect 775 72 776 77
rect 769 71 776 72
rect 985 77 992 78
rect 985 72 986 77
rect 991 72 992 77
rect 985 71 992 72
rect 19 67 26 68
rect 19 62 20 67
rect 25 66 26 67
rect 122 66 126 71
rect 25 62 126 66
rect 235 67 242 68
rect 235 62 236 67
rect 241 66 242 67
rect 338 66 342 71
rect 241 62 342 66
rect 451 67 458 68
rect 451 62 452 67
rect 457 66 458 67
rect 554 66 558 71
rect 457 62 558 66
rect 667 67 674 68
rect 667 62 668 67
rect 673 66 674 67
rect 770 66 774 71
rect 673 62 774 66
rect 883 67 890 68
rect 883 62 884 67
rect 889 66 890 67
rect 986 66 990 71
rect 889 62 990 66
rect 19 61 26 62
rect 235 61 242 62
rect 451 61 458 62
rect 667 61 674 62
rect 883 61 890 62
rect 33 25 62 26
rect 33 23 59 25
rect 249 25 278 26
rect 249 23 275 25
rect 465 25 494 26
rect 465 23 491 25
rect 681 25 710 26
rect 681 23 707 25
rect 897 25 926 26
rect 897 23 923 25
rect 76 19 83 20
rect 76 14 77 19
rect 82 14 83 19
rect 76 10 83 14
rect 292 19 299 20
rect 292 14 293 19
rect 298 14 299 19
rect 127 11 133 12
rect 126 10 127 11
rect 17 7 127 10
rect 17 -15 20 7
rect 126 6 127 7
rect 132 6 133 11
rect 292 10 299 14
rect 508 19 515 20
rect 508 14 509 19
rect 514 14 515 19
rect 343 11 349 12
rect 342 10 343 11
rect 126 5 133 6
rect 233 7 343 10
rect 233 -15 236 7
rect 342 6 343 7
rect 348 6 349 11
rect 508 10 515 14
rect 724 19 731 20
rect 724 14 725 19
rect 730 14 731 19
rect 559 11 565 12
rect 558 10 559 11
rect 342 5 349 6
rect 449 7 559 10
rect 449 -15 452 7
rect 558 6 559 7
rect 564 6 565 11
rect 724 10 731 14
rect 940 19 947 20
rect 940 14 941 19
rect 946 14 947 19
rect 775 11 781 12
rect 774 10 775 11
rect 558 5 565 6
rect 665 7 775 10
rect 665 -15 668 7
rect 774 6 775 7
rect 780 6 781 11
rect 940 10 947 14
rect 991 11 997 12
rect 990 10 991 11
rect 774 5 781 6
rect 881 7 991 10
rect 881 -15 884 7
rect 990 6 991 7
rect 996 6 997 11
rect 990 5 997 6
rect 17 -19 25 -15
rect 233 -19 241 -15
rect 449 -19 457 -15
rect 665 -19 673 -15
rect 881 -19 889 -15
rect 8 -24 15 -23
rect 22 -24 25 -19
rect 8 -29 9 -24
rect 14 -27 25 -24
rect 224 -24 231 -23
rect 238 -24 241 -19
rect 14 -29 15 -27
rect 8 -30 15 -29
rect 224 -29 225 -24
rect 230 -27 241 -24
rect 440 -24 447 -23
rect 454 -24 457 -19
rect 230 -29 231 -27
rect 224 -30 231 -29
rect 440 -29 441 -24
rect 446 -27 457 -24
rect 656 -24 663 -23
rect 670 -24 673 -19
rect 446 -29 447 -27
rect 440 -30 447 -29
rect 656 -29 657 -24
rect 662 -27 673 -24
rect 872 -24 879 -23
rect 886 -24 889 -19
rect 662 -29 663 -27
rect 656 -30 663 -29
rect 872 -29 873 -24
rect 878 -27 889 -24
rect 878 -29 879 -27
rect 872 -30 879 -29
<< labels >>
rlabel metal1 142 10 142 10 1 gnd
rlabel metal1 358 10 358 10 1 gnd
rlabel metal1 574 10 574 10 1 gnd
rlabel metal1 790 10 790 10 1 gnd
rlabel metal1 1006 10 1006 10 1 gnd
rlabel metal1 141 68 141 68 5 vdd
rlabel metal1 357 68 357 68 5 vdd
rlabel metal1 573 68 573 68 5 vdd
rlabel metal1 789 68 789 68 5 vdd
rlabel metal1 1005 68 1005 68 5 vdd
rlabel metal1 109 -8 113 0 1 input_1
port 1 s
rlabel metal1 325 -8 329 0 1 input_2
port 1 s
rlabel metal1 541 -8 545 0 1 input_3
port 1 s
rlabel metal1 757 -8 761 0 1 input_4
port 1 s
rlabel metal1 973 -8 977 0 1 input_5
port 1 s
rlabel metal1 101 -8 105 0 1 input_2
port 2 s
rlabel metal1 317 -8 321 0 1 input_3
port 2 s
rlabel metal1 533 -8 537 0 1 input_4
port 2 s
rlabel metal1 749 -8 753 0 1 input_5
port 2 s
rlabel metal1 965 -8 969 0 1 input_6
port 2 s
rlabel metal1 92 67 101 71 5 ground
port 5 n
rlabel metal1 308 67 317 71 5 ground
port 5 n
rlabel metal1 524 67 533 71 5 ground
port 5 n
rlabel metal1 740 67 749 71 5 ground
port 5 n
rlabel metal1 956 67 965 71 5 ground
port 5 n
rlabel metal1 91 4 100 8 3 power_supply
port 3 w
rlabel metal1 307 4 316 8 3 power_supply
port 3 w
rlabel metal1 523 4 532 8 3 power_supply
port 3 w
rlabel metal1 739 4 748 8 3 power_supply
port 3 w
rlabel metal1 955 4 964 8 3 power_supply
port 3 w
rlabel metal1 117 39 121 43 7 output
port 4 e
rlabel metal1 333 39 337 43 7 output
port 4 e
rlabel metal1 549 39 553 43 7 output
port 4 e
rlabel metal1 765 39 769 43 7 output
port 4 e
rlabel metal1 981 39 985 43 7 output
port 4 e
rlabel metal1 6 64 6 64 5 vdd
rlabel metal1 222 64 222 64 5 vdd
rlabel metal1 438 64 438 64 5 vdd
rlabel metal1 654 64 654 64 5 vdd
rlabel metal1 870 64 870 64 5 vdd
rlabel metal1 22 24 25 26 7 in1
rlabel metal1 238 24 241 26 7 in2
rlabel metal1 454 24 457 26 7 in3
rlabel metal1 670 24 673 26 7 in4
rlabel metal1 886 24 889 26 7 in5
rlabel m2contact 31 6 31 6 1 in1_inv
rlabel m2contact 247 6 247 6 1 in2_inv
rlabel m2contact 463 6 463 6 1 in3_inv
rlabel m2contact 679 6 679 6 1 in4_inv
rlabel m2contact 895 6 895 6 1 in5_inv
rlabel metal3 57 26 57 26 1 in2
rlabel metal3 273 26 273 26 1 in3
rlabel metal3 489 26 489 26 1 in4
rlabel metal3 705 26 705 26 1 in5
rlabel metal3 921 26 921 26 1 in6
<< end >>
