* XOR Gate Layout
.include TSMC_180nm.txt
.param SUPPLY = 1.8
* width is the universal width parameter - 20*LAMBDA
.global gnd vdd
.option scale=0.09u

* SPICE3 file created from XOR2.ext - technology: scmos

M1000 out in2 in1 w_n191_n85# CMOSP w=20 l=2
+  ad=140 pd=54 as=100 ps=50
M1001 in2 in1 out w_n191_n85# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1002 gnd in1 in1_inv Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=100 ps=60
M1003 vdd in1 in1_inv w_n191_n85# CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1004 in2 in1_inv out Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=70 ps=34
M1005 out in2 in1_inv Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0


Vdd vdd gnd 'SUPPLY'
Va in1 gnd pulse 0 1.8 0 0.01ns 0.01ns 10ns 20ns
Vb in2 gnd pulse 0 1.8 0 0.01ns 0.01ns 20ns 40ns

.tran 100p 50n
.ic v(out) = 0

.control
set hcopypscolor = 1
set color0=white
set color1=black

run

set curplottitle="2024102023_XOR"
plot v(in1)+2, v(in2)+4, v(out)
.endc
.end